library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f4edc287",
    12 => x"86c0c64e",
    13 => x"49f4edc2",
    14 => x"48d4dbc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087e5db",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48111e4f",
    50 => x"7808d4ff",
    51 => x"c14866c4",
    52 => x"58a6c888",
    53 => x"ed059870",
    54 => x"1e4f2687",
    55 => x"c348d4ff",
    56 => x"516878ff",
    57 => x"c14866c4",
    58 => x"58a6c888",
    59 => x"eb059870",
    60 => x"1e4f2687",
    61 => x"d4ff1e73",
    62 => x"7bffc34b",
    63 => x"ffc34a6b",
    64 => x"c8496b7b",
    65 => x"c3b17232",
    66 => x"4a6b7bff",
    67 => x"b27131c8",
    68 => x"6b7bffc3",
    69 => x"7232c849",
    70 => x"c44871b1",
    71 => x"264d2687",
    72 => x"264b264c",
    73 => x"5b5e0e4f",
    74 => x"710e5d5c",
    75 => x"4cd4ff4a",
    76 => x"ffc34972",
    77 => x"c27c7199",
    78 => x"05bfd4db",
    79 => x"66d087c8",
    80 => x"d430c948",
    81 => x"66d058a6",
    82 => x"c329d849",
    83 => x"7c7199ff",
    84 => x"d04966d0",
    85 => x"99ffc329",
    86 => x"66d07c71",
    87 => x"c329c849",
    88 => x"7c7199ff",
    89 => x"c34966d0",
    90 => x"7c7199ff",
    91 => x"29d04972",
    92 => x"7199ffc3",
    93 => x"c94b6c7c",
    94 => x"c34dfff0",
    95 => x"d005abff",
    96 => x"7cffc387",
    97 => x"8dc14b6c",
    98 => x"c387c602",
    99 => x"f002abff",
   100 => x"fe487387",
   101 => x"c01e87c7",
   102 => x"48d4ff49",
   103 => x"c178ffc3",
   104 => x"b7c8c381",
   105 => x"87f104a9",
   106 => x"731e4f26",
   107 => x"c487e71e",
   108 => x"c04bdff8",
   109 => x"f0ffc01e",
   110 => x"fd49f7c1",
   111 => x"86c487e7",
   112 => x"c005a8c1",
   113 => x"d4ff87ea",
   114 => x"78ffc348",
   115 => x"c0c0c0c1",
   116 => x"c01ec0c0",
   117 => x"e9c1f0e1",
   118 => x"87c9fd49",
   119 => x"987086c4",
   120 => x"ff87ca05",
   121 => x"ffc348d4",
   122 => x"cb48c178",
   123 => x"87e6fe87",
   124 => x"fe058bc1",
   125 => x"48c087fd",
   126 => x"1e87e6fc",
   127 => x"d4ff1e73",
   128 => x"78ffc348",
   129 => x"1ec04bd3",
   130 => x"c1f0ffc0",
   131 => x"d4fc49c1",
   132 => x"7086c487",
   133 => x"87ca0598",
   134 => x"c348d4ff",
   135 => x"48c178ff",
   136 => x"f1fd87cb",
   137 => x"058bc187",
   138 => x"c087dbff",
   139 => x"87f1fb48",
   140 => x"5c5b5e0e",
   141 => x"4cd4ff0e",
   142 => x"c687dbfd",
   143 => x"e1c01eea",
   144 => x"49c8c1f0",
   145 => x"c487defb",
   146 => x"02a8c186",
   147 => x"eafe87c8",
   148 => x"c148c087",
   149 => x"dafa87e2",
   150 => x"cf497087",
   151 => x"c699ffff",
   152 => x"c802a9ea",
   153 => x"87d3fe87",
   154 => x"cbc148c0",
   155 => x"7cffc387",
   156 => x"fc4bf1c0",
   157 => x"987087f4",
   158 => x"87ebc002",
   159 => x"ffc01ec0",
   160 => x"49fac1f0",
   161 => x"c487defa",
   162 => x"05987086",
   163 => x"ffc387d9",
   164 => x"c3496c7c",
   165 => x"7c7c7cff",
   166 => x"99c0c17c",
   167 => x"c187c402",
   168 => x"c087d548",
   169 => x"c287d148",
   170 => x"87c405ab",
   171 => x"87c848c0",
   172 => x"fe058bc1",
   173 => x"48c087fd",
   174 => x"1e87e4f9",
   175 => x"dbc21e73",
   176 => x"78c148d4",
   177 => x"d0ff4bc7",
   178 => x"fb78c248",
   179 => x"d0ff87c8",
   180 => x"c078c348",
   181 => x"d0e5c01e",
   182 => x"f949c0c1",
   183 => x"86c487c7",
   184 => x"c105a8c1",
   185 => x"abc24b87",
   186 => x"c087c505",
   187 => x"87f9c048",
   188 => x"ff058bc1",
   189 => x"f7fc87d0",
   190 => x"d8dbc287",
   191 => x"05987058",
   192 => x"1ec187cd",
   193 => x"c1f0ffc0",
   194 => x"d8f849d0",
   195 => x"ff86c487",
   196 => x"ffc348d4",
   197 => x"87e0c478",
   198 => x"58dcdbc2",
   199 => x"c248d0ff",
   200 => x"48d4ff78",
   201 => x"c178ffc3",
   202 => x"87f5f748",
   203 => x"5c5b5e0e",
   204 => x"4a710e5d",
   205 => x"ff4dffc3",
   206 => x"7c754cd4",
   207 => x"c448d0ff",
   208 => x"7c7578c3",
   209 => x"ffc01e72",
   210 => x"49d8c1f0",
   211 => x"c487d6f7",
   212 => x"02987086",
   213 => x"48c087c5",
   214 => x"7587f0c0",
   215 => x"7cfec37c",
   216 => x"d41ec0c8",
   217 => x"dcf54966",
   218 => x"7586c487",
   219 => x"757c757c",
   220 => x"e0dad87c",
   221 => x"6c7c754b",
   222 => x"c5059949",
   223 => x"058bc187",
   224 => x"7c7587f3",
   225 => x"c248d0ff",
   226 => x"f648c178",
   227 => x"ff1e87cf",
   228 => x"d0ff4ad4",
   229 => x"78d1c448",
   230 => x"c17affc3",
   231 => x"87f80589",
   232 => x"731e4f26",
   233 => x"c54b711e",
   234 => x"4adfcdee",
   235 => x"c348d4ff",
   236 => x"486878ff",
   237 => x"02a8fec3",
   238 => x"8ac187c5",
   239 => x"7287ed05",
   240 => x"87c5059a",
   241 => x"eac048c0",
   242 => x"029b7387",
   243 => x"66c887cc",
   244 => x"f449731e",
   245 => x"86c487c5",
   246 => x"66c887c6",
   247 => x"87eefe49",
   248 => x"c348d4ff",
   249 => x"737878ff",
   250 => x"87c5059b",
   251 => x"d048d0ff",
   252 => x"f448c178",
   253 => x"731e87eb",
   254 => x"c04a711e",
   255 => x"48d4ff4b",
   256 => x"ff78ffc3",
   257 => x"c3c448d0",
   258 => x"48d4ff78",
   259 => x"7278ffc3",
   260 => x"f0ffc01e",
   261 => x"f449d1c1",
   262 => x"86c487cb",
   263 => x"cd059870",
   264 => x"1ec0c887",
   265 => x"fd4966cc",
   266 => x"86c487f8",
   267 => x"d0ff4b70",
   268 => x"7378c248",
   269 => x"87e9f348",
   270 => x"5c5b5e0e",
   271 => x"1ec00e5d",
   272 => x"c1f0ffc0",
   273 => x"dcf349c9",
   274 => x"c21ed287",
   275 => x"fd49dcdb",
   276 => x"86c887d0",
   277 => x"84c14cc0",
   278 => x"04acb7d2",
   279 => x"dbc287f8",
   280 => x"49bf97dc",
   281 => x"c199c0c3",
   282 => x"c005a9c0",
   283 => x"dbc287e7",
   284 => x"49bf97e3",
   285 => x"dbc231d0",
   286 => x"4abf97e4",
   287 => x"b17232c8",
   288 => x"97e5dbc2",
   289 => x"71b14abf",
   290 => x"ffffcf4c",
   291 => x"84c19cff",
   292 => x"e7c134ca",
   293 => x"e5dbc287",
   294 => x"c149bf97",
   295 => x"c299c631",
   296 => x"bf97e6db",
   297 => x"2ab7c74a",
   298 => x"dbc2b172",
   299 => x"4abf97e1",
   300 => x"c29dcf4d",
   301 => x"bf97e2db",
   302 => x"ca9ac34a",
   303 => x"e3dbc232",
   304 => x"c24bbf97",
   305 => x"c2b27333",
   306 => x"bf97e4db",
   307 => x"9bc0c34b",
   308 => x"732bb7c6",
   309 => x"c181c2b2",
   310 => x"70307148",
   311 => x"7548c149",
   312 => x"724d7030",
   313 => x"7184c14c",
   314 => x"b7c0c894",
   315 => x"87cc06ad",
   316 => x"2db734c1",
   317 => x"adb7c0c8",
   318 => x"87f4ff01",
   319 => x"dcf04874",
   320 => x"5b5e0e87",
   321 => x"f80e5d5c",
   322 => x"c2e4c286",
   323 => x"c278c048",
   324 => x"c01efadb",
   325 => x"87defb49",
   326 => x"987086c4",
   327 => x"c087c505",
   328 => x"87cec948",
   329 => x"7ec14dc0",
   330 => x"bfcbf2c0",
   331 => x"f0dcc249",
   332 => x"4bc8714a",
   333 => x"7087f3ec",
   334 => x"87c20598",
   335 => x"f2c07ec0",
   336 => x"c249bfc7",
   337 => x"714accdd",
   338 => x"ddec4bc8",
   339 => x"05987087",
   340 => x"7ec087c2",
   341 => x"fdc0026e",
   342 => x"c0e3c287",
   343 => x"e3c24dbf",
   344 => x"7ebf9ff8",
   345 => x"ead6c548",
   346 => x"87c705a8",
   347 => x"bfc0e3c2",
   348 => x"6e87ce4d",
   349 => x"d5e9ca48",
   350 => x"87c502a8",
   351 => x"f1c748c0",
   352 => x"fadbc287",
   353 => x"f949751e",
   354 => x"86c487ec",
   355 => x"c5059870",
   356 => x"c748c087",
   357 => x"f2c087dc",
   358 => x"c249bfc7",
   359 => x"714accdd",
   360 => x"c5eb4bc8",
   361 => x"05987087",
   362 => x"e4c287c8",
   363 => x"78c148c2",
   364 => x"f2c087da",
   365 => x"c249bfcb",
   366 => x"714af0dc",
   367 => x"e9ea4bc8",
   368 => x"02987087",
   369 => x"c087c5c0",
   370 => x"87e6c648",
   371 => x"97f8e3c2",
   372 => x"d5c149bf",
   373 => x"cdc005a9",
   374 => x"f9e3c287",
   375 => x"c249bf97",
   376 => x"c002a9ea",
   377 => x"48c087c5",
   378 => x"c287c7c6",
   379 => x"bf97fadb",
   380 => x"e9c3487e",
   381 => x"cec002a8",
   382 => x"c3486e87",
   383 => x"c002a8eb",
   384 => x"48c087c5",
   385 => x"c287ebc5",
   386 => x"bf97c5dc",
   387 => x"c0059949",
   388 => x"dcc287cc",
   389 => x"49bf97c6",
   390 => x"c002a9c2",
   391 => x"48c087c5",
   392 => x"c287cfc5",
   393 => x"bf97c7dc",
   394 => x"fee3c248",
   395 => x"484c7058",
   396 => x"e4c288c1",
   397 => x"dcc258c2",
   398 => x"49bf97c8",
   399 => x"dcc28175",
   400 => x"4abf97c9",
   401 => x"a17232c8",
   402 => x"cfe8c27e",
   403 => x"c2786e48",
   404 => x"bf97cadc",
   405 => x"58a6c848",
   406 => x"bfc2e4c2",
   407 => x"87d4c202",
   408 => x"bfc7f2c0",
   409 => x"ccddc249",
   410 => x"4bc8714a",
   411 => x"7087fbe7",
   412 => x"c5c00298",
   413 => x"c348c087",
   414 => x"e3c287f8",
   415 => x"c24cbffa",
   416 => x"c25ce3e8",
   417 => x"bf97dfdc",
   418 => x"c231c849",
   419 => x"bf97dedc",
   420 => x"c249a14a",
   421 => x"bf97e0dc",
   422 => x"7232d04a",
   423 => x"dcc249a1",
   424 => x"4abf97e1",
   425 => x"a17232d8",
   426 => x"9166c449",
   427 => x"bfcfe8c2",
   428 => x"d7e8c281",
   429 => x"e7dcc259",
   430 => x"c84abf97",
   431 => x"e6dcc232",
   432 => x"a24bbf97",
   433 => x"e8dcc24a",
   434 => x"d04bbf97",
   435 => x"4aa27333",
   436 => x"97e9dcc2",
   437 => x"9bcf4bbf",
   438 => x"a27333d8",
   439 => x"dbe8c24a",
   440 => x"d7e8c25a",
   441 => x"8ac24abf",
   442 => x"e8c29274",
   443 => x"a17248db",
   444 => x"87cac178",
   445 => x"97ccdcc2",
   446 => x"31c849bf",
   447 => x"97cbdcc2",
   448 => x"49a14abf",
   449 => x"59cae4c2",
   450 => x"bfc6e4c2",
   451 => x"c731c549",
   452 => x"29c981ff",
   453 => x"59e3e8c2",
   454 => x"97d1dcc2",
   455 => x"32c84abf",
   456 => x"97d0dcc2",
   457 => x"4aa24bbf",
   458 => x"6e9266c4",
   459 => x"dfe8c282",
   460 => x"d7e8c25a",
   461 => x"c278c048",
   462 => x"7248d3e8",
   463 => x"e8c278a1",
   464 => x"e8c248e3",
   465 => x"c278bfd7",
   466 => x"c248e7e8",
   467 => x"78bfdbe8",
   468 => x"bfc2e4c2",
   469 => x"87c9c002",
   470 => x"30c44874",
   471 => x"c9c07e70",
   472 => x"dfe8c287",
   473 => x"30c448bf",
   474 => x"e4c27e70",
   475 => x"786e48c6",
   476 => x"8ef848c1",
   477 => x"4c264d26",
   478 => x"4f264b26",
   479 => x"5c5b5e0e",
   480 => x"4a710e5d",
   481 => x"bfc2e4c2",
   482 => x"7287cb02",
   483 => x"722bc74b",
   484 => x"9cffc14c",
   485 => x"4b7287c9",
   486 => x"4c722bc8",
   487 => x"c29cffc3",
   488 => x"83bfcfe8",
   489 => x"bfc3f2c0",
   490 => x"87d902ab",
   491 => x"5bc7f2c0",
   492 => x"1efadbc2",
   493 => x"fdf04973",
   494 => x"7086c487",
   495 => x"87c50598",
   496 => x"e6c048c0",
   497 => x"c2e4c287",
   498 => x"87d202bf",
   499 => x"91c44974",
   500 => x"81fadbc2",
   501 => x"ffcf4d69",
   502 => x"9dffffff",
   503 => x"497487cb",
   504 => x"dbc291c2",
   505 => x"699f81fa",
   506 => x"fe48754d",
   507 => x"5e0e87c6",
   508 => x"0e5d5c5b",
   509 => x"c04d711e",
   510 => x"ca49c11e",
   511 => x"86c487ee",
   512 => x"029c4c70",
   513 => x"c287c0c1",
   514 => x"754acae4",
   515 => x"87ffe049",
   516 => x"c0029870",
   517 => x"4a7487f1",
   518 => x"4bcb4975",
   519 => x"7087e5e1",
   520 => x"e2c00298",
   521 => x"741ec087",
   522 => x"87c7029c",
   523 => x"c048a6c4",
   524 => x"c487c578",
   525 => x"78c148a6",
   526 => x"c94966c4",
   527 => x"86c487ee",
   528 => x"059c4c70",
   529 => x"7487c0ff",
   530 => x"e7fc2648",
   531 => x"5b5e0e87",
   532 => x"1e0e5d5c",
   533 => x"059b4b71",
   534 => x"48c087c5",
   535 => x"c887e5c1",
   536 => x"7dc04da3",
   537 => x"c70266d4",
   538 => x"9766d487",
   539 => x"87c505bf",
   540 => x"cfc148c0",
   541 => x"4966d487",
   542 => x"7087f3fd",
   543 => x"c1029c4c",
   544 => x"a4dc87c0",
   545 => x"da7d6949",
   546 => x"a3c449a4",
   547 => x"7a699f4a",
   548 => x"bfc2e4c2",
   549 => x"d487d202",
   550 => x"699f49a4",
   551 => x"ffffc049",
   552 => x"d0487199",
   553 => x"c27e7030",
   554 => x"6e7ec087",
   555 => x"806a4849",
   556 => x"7bc07a70",
   557 => x"6a49a3cc",
   558 => x"49a3d079",
   559 => x"487479c0",
   560 => x"48c087c2",
   561 => x"87ecfa26",
   562 => x"5c5b5e0e",
   563 => x"4c710e5d",
   564 => x"48c3f2c0",
   565 => x"9c7478ff",
   566 => x"87cac102",
   567 => x"6949a4c8",
   568 => x"87c2c102",
   569 => x"6c4a66d0",
   570 => x"a6d48249",
   571 => x"4d66d05a",
   572 => x"fee3c2b9",
   573 => x"baff4abf",
   574 => x"99719972",
   575 => x"87e4c002",
   576 => x"6b4ba4c4",
   577 => x"87f4f949",
   578 => x"e3c27b70",
   579 => x"6c49bffa",
   580 => x"757c7181",
   581 => x"fee3c2b9",
   582 => x"baff4abf",
   583 => x"99719972",
   584 => x"87dcff05",
   585 => x"cbf97c75",
   586 => x"1e731e87",
   587 => x"029b4b71",
   588 => x"a3c887c7",
   589 => x"c5056949",
   590 => x"c048c087",
   591 => x"e8c287eb",
   592 => x"c44abfd3",
   593 => x"496949a3",
   594 => x"e3c289c2",
   595 => x"7191bffa",
   596 => x"e3c24aa2",
   597 => x"6b49bffe",
   598 => x"4aa27199",
   599 => x"721e66c8",
   600 => x"87d2ea49",
   601 => x"497086c4",
   602 => x"87ccf848",
   603 => x"711e731e",
   604 => x"c7029b4b",
   605 => x"49a3c887",
   606 => x"87c50569",
   607 => x"ebc048c0",
   608 => x"d3e8c287",
   609 => x"a3c44abf",
   610 => x"c2496949",
   611 => x"fae3c289",
   612 => x"a27191bf",
   613 => x"fee3c24a",
   614 => x"996b49bf",
   615 => x"c84aa271",
   616 => x"49721e66",
   617 => x"c487c5e6",
   618 => x"48497086",
   619 => x"0e87c9f7",
   620 => x"5d5c5b5e",
   621 => x"4b711e0e",
   622 => x"c94c66d4",
   623 => x"029b732c",
   624 => x"c887cfc1",
   625 => x"026949a3",
   626 => x"d087c7c1",
   627 => x"66d44da3",
   628 => x"fee3c27d",
   629 => x"b9ff49bf",
   630 => x"7e994a6b",
   631 => x"cd03ac71",
   632 => x"7d7bc087",
   633 => x"c44aa3cc",
   634 => x"796a49a3",
   635 => x"8c7287c2",
   636 => x"dd029c74",
   637 => x"731e4987",
   638 => x"87ccfb49",
   639 => x"66d486c4",
   640 => x"99ffc749",
   641 => x"c287cb02",
   642 => x"731efadb",
   643 => x"87d9fc49",
   644 => x"f52686c4",
   645 => x"731e87de",
   646 => x"9b4b711e",
   647 => x"87e4c002",
   648 => x"5be7e8c2",
   649 => x"8ac24a73",
   650 => x"bffae3c2",
   651 => x"e8c29249",
   652 => x"7248bfd3",
   653 => x"ebe8c280",
   654 => x"c4487158",
   655 => x"cae4c230",
   656 => x"87edc058",
   657 => x"48e3e8c2",
   658 => x"bfd7e8c2",
   659 => x"e7e8c278",
   660 => x"dbe8c248",
   661 => x"e4c278bf",
   662 => x"c902bfc2",
   663 => x"fae3c287",
   664 => x"31c449bf",
   665 => x"e8c287c7",
   666 => x"c449bfdf",
   667 => x"cae4c231",
   668 => x"87c4f459",
   669 => x"5c5b5e0e",
   670 => x"c04a710e",
   671 => x"029a724b",
   672 => x"da87e1c0",
   673 => x"699f49a2",
   674 => x"c2e4c24b",
   675 => x"87cf02bf",
   676 => x"9f49a2d4",
   677 => x"c04c4969",
   678 => x"d09cffff",
   679 => x"c087c234",
   680 => x"b349744c",
   681 => x"edfd4973",
   682 => x"87caf387",
   683 => x"5c5b5e0e",
   684 => x"86f40e5d",
   685 => x"7ec04a71",
   686 => x"d8029a72",
   687 => x"f6dbc287",
   688 => x"c278c048",
   689 => x"c248eedb",
   690 => x"78bfe7e8",
   691 => x"48f2dbc2",
   692 => x"bfe3e8c2",
   693 => x"d7e4c278",
   694 => x"c250c048",
   695 => x"49bfc6e4",
   696 => x"bff6dbc2",
   697 => x"03aa714a",
   698 => x"7287ffc3",
   699 => x"0599cf49",
   700 => x"c287e0c0",
   701 => x"c21efadb",
   702 => x"49bfeedb",
   703 => x"48eedbc2",
   704 => x"7178a1c1",
   705 => x"c487efe3",
   706 => x"fff1c086",
   707 => x"fadbc248",
   708 => x"c087cc78",
   709 => x"48bffff1",
   710 => x"c080e0c0",
   711 => x"c258c3f2",
   712 => x"48bff6db",
   713 => x"dbc280c1",
   714 => x"7f2758fa",
   715 => x"bf00000c",
   716 => x"9d4dbf97",
   717 => x"87e2c202",
   718 => x"02ade5c3",
   719 => x"c087dbc2",
   720 => x"4bbffff1",
   721 => x"1149a3cb",
   722 => x"05accf4c",
   723 => x"7587d2c1",
   724 => x"c199df49",
   725 => x"c291cd89",
   726 => x"c181cae4",
   727 => x"51124aa3",
   728 => x"124aa3c3",
   729 => x"4aa3c551",
   730 => x"a3c75112",
   731 => x"c951124a",
   732 => x"51124aa3",
   733 => x"124aa3ce",
   734 => x"4aa3d051",
   735 => x"a3d25112",
   736 => x"d451124a",
   737 => x"51124aa3",
   738 => x"124aa3d6",
   739 => x"4aa3d851",
   740 => x"a3dc5112",
   741 => x"de51124a",
   742 => x"51124aa3",
   743 => x"f9c07ec1",
   744 => x"c8497487",
   745 => x"eac00599",
   746 => x"d0497487",
   747 => x"87d00599",
   748 => x"c00266dc",
   749 => x"497387ca",
   750 => x"700f66dc",
   751 => x"87d30298",
   752 => x"c6c0056e",
   753 => x"cae4c287",
   754 => x"c050c048",
   755 => x"48bffff1",
   756 => x"c287e7c2",
   757 => x"c048d7e4",
   758 => x"e4c27e50",
   759 => x"c249bfc6",
   760 => x"4abff6db",
   761 => x"fc04aa71",
   762 => x"e8c287c1",
   763 => x"c005bfe7",
   764 => x"e4c287c8",
   765 => x"c102bfc2",
   766 => x"f2c087fe",
   767 => x"78ff48c3",
   768 => x"bff2dbc2",
   769 => x"87f4ed49",
   770 => x"dbc24970",
   771 => x"a6c459f6",
   772 => x"f2dbc248",
   773 => x"e4c278bf",
   774 => x"c002bfc2",
   775 => x"66c487d8",
   776 => x"ffffcf49",
   777 => x"a999f8ff",
   778 => x"87c5c002",
   779 => x"e1c04dc0",
   780 => x"c04dc187",
   781 => x"66c487dc",
   782 => x"f8ffcf49",
   783 => x"c002a999",
   784 => x"a6c887c8",
   785 => x"c078c048",
   786 => x"a6c887c5",
   787 => x"c878c148",
   788 => x"9d754d66",
   789 => x"87e0c005",
   790 => x"c24966c4",
   791 => x"fae3c289",
   792 => x"c2914abf",
   793 => x"4abfd3e8",
   794 => x"48eedbc2",
   795 => x"c278a172",
   796 => x"c048f6db",
   797 => x"87e3f978",
   798 => x"8ef448c0",
   799 => x"0087f5eb",
   800 => x"ff000000",
   801 => x"8fffffff",
   802 => x"9800000c",
   803 => x"4600000c",
   804 => x"32335441",
   805 => x"00202020",
   806 => x"31544146",
   807 => x"20202036",
   808 => x"d4ff1e00",
   809 => x"78ffc348",
   810 => x"4f264868",
   811 => x"48d4ff1e",
   812 => x"ff78ffc3",
   813 => x"e1c848d0",
   814 => x"48d4ff78",
   815 => x"e8c278d4",
   816 => x"d4ff48eb",
   817 => x"4f2650bf",
   818 => x"48d0ff1e",
   819 => x"2678e0c0",
   820 => x"ccff1e4f",
   821 => x"99497087",
   822 => x"c087c602",
   823 => x"f105a9fb",
   824 => x"26487187",
   825 => x"5b5e0e4f",
   826 => x"4b710e5c",
   827 => x"f0fe4cc0",
   828 => x"99497087",
   829 => x"87f9c002",
   830 => x"02a9ecc0",
   831 => x"c087f2c0",
   832 => x"c002a9fb",
   833 => x"66cc87eb",
   834 => x"c703acb7",
   835 => x"0266d087",
   836 => x"537187c2",
   837 => x"c2029971",
   838 => x"fe84c187",
   839 => x"497087c3",
   840 => x"87cd0299",
   841 => x"02a9ecc0",
   842 => x"fbc087c7",
   843 => x"d5ff05a9",
   844 => x"0266d087",
   845 => x"97c087c3",
   846 => x"a9ecc07b",
   847 => x"7487c405",
   848 => x"7487c54a",
   849 => x"8a0ac04a",
   850 => x"87c24872",
   851 => x"4c264d26",
   852 => x"4f264b26",
   853 => x"87c9fd1e",
   854 => x"f0c04970",
   855 => x"ca04a9b7",
   856 => x"b7f9c087",
   857 => x"87c301a9",
   858 => x"c189f0c0",
   859 => x"04a9b7c1",
   860 => x"dac187ca",
   861 => x"c301a9b7",
   862 => x"89f7c087",
   863 => x"4f264871",
   864 => x"5c5b5e0e",
   865 => x"ff4a710e",
   866 => x"49724cd4",
   867 => x"7087eac0",
   868 => x"c2029b4b",
   869 => x"ff8bc187",
   870 => x"c5c848d0",
   871 => x"7cd5c178",
   872 => x"31c64973",
   873 => x"97e4dac2",
   874 => x"71484abf",
   875 => x"ff7c70b0",
   876 => x"78c448d0",
   877 => x"d5fe4873",
   878 => x"5b5e0e87",
   879 => x"f80e5d5c",
   880 => x"c04c7186",
   881 => x"87e4fb7e",
   882 => x"f9c04bc0",
   883 => x"49bf97e6",
   884 => x"cf04a9c0",
   885 => x"87f9fb87",
   886 => x"f9c083c1",
   887 => x"49bf97e6",
   888 => x"87f106ab",
   889 => x"97e6f9c0",
   890 => x"87cf02bf",
   891 => x"7087f2fa",
   892 => x"c6029949",
   893 => x"a9ecc087",
   894 => x"c087f105",
   895 => x"87e1fa4b",
   896 => x"dcfa4d70",
   897 => x"58a6c887",
   898 => x"7087d6fa",
   899 => x"c883c14a",
   900 => x"699749a4",
   901 => x"c702ad49",
   902 => x"adffc087",
   903 => x"87e7c005",
   904 => x"9749a4c9",
   905 => x"66c44969",
   906 => x"87c702a9",
   907 => x"a8ffc048",
   908 => x"ca87d405",
   909 => x"699749a4",
   910 => x"c602aa49",
   911 => x"aaffc087",
   912 => x"c187c405",
   913 => x"c087d07e",
   914 => x"c602adec",
   915 => x"adfbc087",
   916 => x"c087c405",
   917 => x"6e7ec14b",
   918 => x"87e1fe02",
   919 => x"7387e9f9",
   920 => x"fb8ef848",
   921 => x"0e0087e6",
   922 => x"5d5c5b5e",
   923 => x"4b711e0e",
   924 => x"ab4d4cc0",
   925 => x"87e8c004",
   926 => x"1ef9f6c0",
   927 => x"c4029d75",
   928 => x"c24ac087",
   929 => x"724ac187",
   930 => x"87e0f049",
   931 => x"7e7086c4",
   932 => x"056e84c1",
   933 => x"4c7387c2",
   934 => x"ac7385c1",
   935 => x"87d8ff06",
   936 => x"2626486e",
   937 => x"264c264d",
   938 => x"0e4f264b",
   939 => x"5d5c5b5e",
   940 => x"4c711e0e",
   941 => x"c291de49",
   942 => x"714dc5e9",
   943 => x"026d9785",
   944 => x"c287ddc1",
   945 => x"4abff0e8",
   946 => x"49728274",
   947 => x"7087d8fe",
   948 => x"c0026e7e",
   949 => x"e8c287f3",
   950 => x"4a6e4bf8",
   951 => x"c7ff49cb",
   952 => x"4b7487c6",
   953 => x"ddc193cb",
   954 => x"83c483d4",
   955 => x"7be4fcc0",
   956 => x"c3c14974",
   957 => x"7b7587c5",
   958 => x"97c4e9c2",
   959 => x"c21e49bf",
   960 => x"c149f8e8",
   961 => x"c487dfdd",
   962 => x"c1497486",
   963 => x"c087ecc2",
   964 => x"cbc4c149",
   965 => x"ece8c287",
   966 => x"c178c048",
   967 => x"87cbdd49",
   968 => x"87fffd26",
   969 => x"64616f4c",
   970 => x"2e676e69",
   971 => x"0e002e2e",
   972 => x"0e5c5b5e",
   973 => x"c24a4b71",
   974 => x"82bff0e8",
   975 => x"e6fc4972",
   976 => x"9c4c7087",
   977 => x"4987c402",
   978 => x"c287e9ec",
   979 => x"c048f0e8",
   980 => x"dc49c178",
   981 => x"ccfd87d5",
   982 => x"5b5e0e87",
   983 => x"f40e5d5c",
   984 => x"fadbc286",
   985 => x"c44cc04d",
   986 => x"78c048a6",
   987 => x"bff0e8c2",
   988 => x"06a9c049",
   989 => x"c287c1c1",
   990 => x"9848fadb",
   991 => x"87f8c002",
   992 => x"1ef9f6c0",
   993 => x"c70266c8",
   994 => x"48a6c487",
   995 => x"87c578c0",
   996 => x"c148a6c4",
   997 => x"4966c478",
   998 => x"c487d1ec",
   999 => x"c14d7086",
  1000 => x"4866c484",
  1001 => x"a6c880c1",
  1002 => x"f0e8c258",
  1003 => x"03ac49bf",
  1004 => x"9d7587c6",
  1005 => x"87c8ff05",
  1006 => x"9d754cc0",
  1007 => x"87e0c302",
  1008 => x"1ef9f6c0",
  1009 => x"c70266c8",
  1010 => x"48a6cc87",
  1011 => x"87c578c0",
  1012 => x"c148a6cc",
  1013 => x"4966cc78",
  1014 => x"c487d1eb",
  1015 => x"6e7e7086",
  1016 => x"87e9c202",
  1017 => x"81cb496e",
  1018 => x"d0496997",
  1019 => x"d6c10299",
  1020 => x"effcc087",
  1021 => x"cb49744a",
  1022 => x"d4ddc191",
  1023 => x"c8797281",
  1024 => x"51ffc381",
  1025 => x"91de4974",
  1026 => x"4dc5e9c2",
  1027 => x"c1c28571",
  1028 => x"a5c17d97",
  1029 => x"51e0c049",
  1030 => x"97cae4c2",
  1031 => x"87d202bf",
  1032 => x"a5c284c1",
  1033 => x"cae4c24b",
  1034 => x"ff49db4a",
  1035 => x"c187f9c1",
  1036 => x"a5cd87db",
  1037 => x"c151c049",
  1038 => x"4ba5c284",
  1039 => x"49cb4a6e",
  1040 => x"87e4c1ff",
  1041 => x"c087c6c1",
  1042 => x"744aebfa",
  1043 => x"c191cb49",
  1044 => x"7281d4dd",
  1045 => x"cae4c279",
  1046 => x"d802bf97",
  1047 => x"de497487",
  1048 => x"c284c191",
  1049 => x"714bc5e9",
  1050 => x"cae4c283",
  1051 => x"ff49dd4a",
  1052 => x"d887f5c0",
  1053 => x"de4b7487",
  1054 => x"c5e9c293",
  1055 => x"49a3cb83",
  1056 => x"84c151c0",
  1057 => x"cb4a6e73",
  1058 => x"dbc0ff49",
  1059 => x"4866c487",
  1060 => x"a6c880c1",
  1061 => x"03acc758",
  1062 => x"6e87c5c0",
  1063 => x"87e0fc05",
  1064 => x"8ef44874",
  1065 => x"1e87fcf7",
  1066 => x"4b711e73",
  1067 => x"c191cb49",
  1068 => x"c881d4dd",
  1069 => x"dac24aa1",
  1070 => x"501248e4",
  1071 => x"c04aa1c9",
  1072 => x"1248e6f9",
  1073 => x"c281ca50",
  1074 => x"1148c4e9",
  1075 => x"c4e9c250",
  1076 => x"1e49bf97",
  1077 => x"d6c149c0",
  1078 => x"e8c287cc",
  1079 => x"78de48ec",
  1080 => x"c6d649c1",
  1081 => x"fef62687",
  1082 => x"4a711e87",
  1083 => x"c191cb49",
  1084 => x"c881d4dd",
  1085 => x"c2481181",
  1086 => x"c258f0e8",
  1087 => x"c048f0e8",
  1088 => x"d549c178",
  1089 => x"4f2687e5",
  1090 => x"c049c01e",
  1091 => x"2687d1fc",
  1092 => x"99711e4f",
  1093 => x"c187d202",
  1094 => x"c048e9de",
  1095 => x"c180f750",
  1096 => x"c140e9c3",
  1097 => x"ce78cddd",
  1098 => x"e5dec187",
  1099 => x"c6ddc148",
  1100 => x"c180fc78",
  1101 => x"2678c8c4",
  1102 => x"5b5e0e4f",
  1103 => x"4c710e5c",
  1104 => x"c192cb4a",
  1105 => x"c882d4dd",
  1106 => x"a2c949a2",
  1107 => x"4b6b974b",
  1108 => x"4969971e",
  1109 => x"1282ca1e",
  1110 => x"cce7c049",
  1111 => x"d449c087",
  1112 => x"497487c9",
  1113 => x"87d3f9c0",
  1114 => x"f8f48ef8",
  1115 => x"1e731e87",
  1116 => x"ff494b71",
  1117 => x"497387c3",
  1118 => x"f487fefe",
  1119 => x"731e87e9",
  1120 => x"c64b711e",
  1121 => x"db024aa3",
  1122 => x"028ac187",
  1123 => x"028a87d6",
  1124 => x"8a87dac1",
  1125 => x"87fcc002",
  1126 => x"e1c0028a",
  1127 => x"cb028a87",
  1128 => x"87dbc187",
  1129 => x"c0fd49c7",
  1130 => x"87dec187",
  1131 => x"bff0e8c2",
  1132 => x"87cbc102",
  1133 => x"c288c148",
  1134 => x"c158f4e8",
  1135 => x"e8c287c1",
  1136 => x"c002bff4",
  1137 => x"e8c287f9",
  1138 => x"c148bff0",
  1139 => x"f4e8c280",
  1140 => x"87ebc058",
  1141 => x"bff0e8c2",
  1142 => x"c289c649",
  1143 => x"c059f4e8",
  1144 => x"da03a9b7",
  1145 => x"f0e8c287",
  1146 => x"d278c048",
  1147 => x"f4e8c287",
  1148 => x"87cb02bf",
  1149 => x"bff0e8c2",
  1150 => x"c280c648",
  1151 => x"c058f4e8",
  1152 => x"87e7d149",
  1153 => x"f6c04973",
  1154 => x"daf287f1",
  1155 => x"5b5e0e87",
  1156 => x"4c710e5c",
  1157 => x"741e66cc",
  1158 => x"c193cb4b",
  1159 => x"c483d4dd",
  1160 => x"496a4aa3",
  1161 => x"87d0fafe",
  1162 => x"7be7c2c1",
  1163 => x"d449a3c8",
  1164 => x"a3c95166",
  1165 => x"5166d849",
  1166 => x"dc49a3ca",
  1167 => x"f1265166",
  1168 => x"5e0e87e3",
  1169 => x"0e5d5c5b",
  1170 => x"d886d0ff",
  1171 => x"a6c459a6",
  1172 => x"c478c048",
  1173 => x"66c4c180",
  1174 => x"c180c478",
  1175 => x"c180c478",
  1176 => x"f4e8c278",
  1177 => x"c278c148",
  1178 => x"48bfece8",
  1179 => x"cb05a8de",
  1180 => x"87e5f387",
  1181 => x"a6c84970",
  1182 => x"87f8ce59",
  1183 => x"e987ede8",
  1184 => x"dce887cf",
  1185 => x"c04c7087",
  1186 => x"c102acfb",
  1187 => x"66d487d0",
  1188 => x"87c2c105",
  1189 => x"c11e1ec0",
  1190 => x"c7dfc11e",
  1191 => x"fd49c01e",
  1192 => x"d0c187eb",
  1193 => x"82c44a66",
  1194 => x"81c7496a",
  1195 => x"1ec15174",
  1196 => x"496a1ed8",
  1197 => x"ece881c8",
  1198 => x"c186d887",
  1199 => x"c04866c4",
  1200 => x"87c701a8",
  1201 => x"c148a6c4",
  1202 => x"c187ce78",
  1203 => x"c14866c4",
  1204 => x"58a6cc88",
  1205 => x"f8e787c3",
  1206 => x"48a6cc87",
  1207 => x"9c7478c2",
  1208 => x"87cccd02",
  1209 => x"c14866c4",
  1210 => x"03a866c8",
  1211 => x"d887c1cd",
  1212 => x"78c048a6",
  1213 => x"7087eae6",
  1214 => x"acd0c14c",
  1215 => x"87d6c205",
  1216 => x"e97e66d8",
  1217 => x"497087ce",
  1218 => x"e659a6dc",
  1219 => x"4c7087d3",
  1220 => x"05acecc0",
  1221 => x"c487eac1",
  1222 => x"91cb4966",
  1223 => x"8166c0c1",
  1224 => x"6a4aa1c4",
  1225 => x"4aa1c84d",
  1226 => x"c15266d8",
  1227 => x"e579e9c3",
  1228 => x"4c7087ef",
  1229 => x"87d8029c",
  1230 => x"02acfbc0",
  1231 => x"557487d2",
  1232 => x"7087dee5",
  1233 => x"c7029c4c",
  1234 => x"acfbc087",
  1235 => x"87eeff05",
  1236 => x"c255e0c0",
  1237 => x"97c055c1",
  1238 => x"4966d47d",
  1239 => x"db05a96e",
  1240 => x"4866c487",
  1241 => x"04a866c8",
  1242 => x"66c487ca",
  1243 => x"c880c148",
  1244 => x"87c858a6",
  1245 => x"c14866c8",
  1246 => x"58a6cc88",
  1247 => x"7087e2e4",
  1248 => x"acd0c14c",
  1249 => x"d087c805",
  1250 => x"80c14866",
  1251 => x"c158a6d4",
  1252 => x"fd02acd0",
  1253 => x"a6dc87ea",
  1254 => x"7866d448",
  1255 => x"dc4866d8",
  1256 => x"c905a866",
  1257 => x"e0c087dc",
  1258 => x"f0c048a6",
  1259 => x"cc80c478",
  1260 => x"80c47866",
  1261 => x"747e78c0",
  1262 => x"88fbc048",
  1263 => x"58a6f0c0",
  1264 => x"c8029870",
  1265 => x"cb4887d7",
  1266 => x"a6f0c088",
  1267 => x"02987058",
  1268 => x"4887e9c0",
  1269 => x"f0c088c9",
  1270 => x"987058a6",
  1271 => x"87e1c302",
  1272 => x"c088c448",
  1273 => x"7058a6f0",
  1274 => x"87d60298",
  1275 => x"c088c148",
  1276 => x"7058a6f0",
  1277 => x"c8c30298",
  1278 => x"87dbc787",
  1279 => x"48a6e0c0",
  1280 => x"66cc78c0",
  1281 => x"d080c148",
  1282 => x"d4e258a6",
  1283 => x"c04c7087",
  1284 => x"d502acec",
  1285 => x"66e0c087",
  1286 => x"c087c602",
  1287 => x"c95ca6e4",
  1288 => x"c0487487",
  1289 => x"e8c088f0",
  1290 => x"ecc058a6",
  1291 => x"87cc02ac",
  1292 => x"7087eee1",
  1293 => x"acecc04c",
  1294 => x"87f4ff05",
  1295 => x"1e66e0c0",
  1296 => x"1e4966d4",
  1297 => x"1e66ecc0",
  1298 => x"1ec7dfc1",
  1299 => x"f64966d4",
  1300 => x"1ec087fb",
  1301 => x"66dc1eca",
  1302 => x"c191cb49",
  1303 => x"d88166d8",
  1304 => x"a1c448a6",
  1305 => x"bf66d878",
  1306 => x"87f9e149",
  1307 => x"b7c086d8",
  1308 => x"c7c106a8",
  1309 => x"de1ec187",
  1310 => x"bf66c81e",
  1311 => x"87e5e149",
  1312 => x"497086c8",
  1313 => x"8808c048",
  1314 => x"58a6e4c0",
  1315 => x"06a8b7c0",
  1316 => x"c087e9c0",
  1317 => x"dd4866e0",
  1318 => x"df03a8b7",
  1319 => x"49bf6e87",
  1320 => x"8166e0c0",
  1321 => x"6651e0c0",
  1322 => x"6e81c149",
  1323 => x"c1c281bf",
  1324 => x"66e0c051",
  1325 => x"6e81c249",
  1326 => x"51c081bf",
  1327 => x"dcc47ec1",
  1328 => x"87d0e287",
  1329 => x"58a6e4c0",
  1330 => x"c087c9e2",
  1331 => x"c058a6e8",
  1332 => x"c005a8ec",
  1333 => x"e4c087cb",
  1334 => x"e0c048a6",
  1335 => x"c4c07866",
  1336 => x"fcdeff87",
  1337 => x"4966c487",
  1338 => x"c0c191cb",
  1339 => x"80714866",
  1340 => x"4a6e7e70",
  1341 => x"496e82c8",
  1342 => x"e0c081ca",
  1343 => x"e4c05166",
  1344 => x"81c14966",
  1345 => x"8966e0c0",
  1346 => x"307148c1",
  1347 => x"89c14970",
  1348 => x"c27a9771",
  1349 => x"49bfe1ec",
  1350 => x"2966e0c0",
  1351 => x"484a6a97",
  1352 => x"f0c09871",
  1353 => x"496e58a6",
  1354 => x"4d6981c4",
  1355 => x"d84866dc",
  1356 => x"c002a866",
  1357 => x"a6d887c8",
  1358 => x"c078c048",
  1359 => x"a6d887c5",
  1360 => x"d878c148",
  1361 => x"e0c01e66",
  1362 => x"ff49751e",
  1363 => x"c887d6de",
  1364 => x"c04c7086",
  1365 => x"c106acb7",
  1366 => x"857487d4",
  1367 => x"7449e0c0",
  1368 => x"c14b7589",
  1369 => x"714ae8d9",
  1370 => x"87fcecfe",
  1371 => x"e8c085c2",
  1372 => x"80c14866",
  1373 => x"58a6ecc0",
  1374 => x"4966ecc0",
  1375 => x"a97081c1",
  1376 => x"87c8c002",
  1377 => x"c048a6d8",
  1378 => x"87c5c078",
  1379 => x"c148a6d8",
  1380 => x"1e66d878",
  1381 => x"c049a4c2",
  1382 => x"887148e0",
  1383 => x"751e4970",
  1384 => x"c0ddff49",
  1385 => x"c086c887",
  1386 => x"ff01a8b7",
  1387 => x"e8c087c0",
  1388 => x"d1c00266",
  1389 => x"c9496e87",
  1390 => x"66e8c081",
  1391 => x"c1486e51",
  1392 => x"c078f9c4",
  1393 => x"496e87cc",
  1394 => x"51c281c9",
  1395 => x"c5c1486e",
  1396 => x"7ec178ed",
  1397 => x"ff87c6c0",
  1398 => x"7087f6db",
  1399 => x"c0026e4c",
  1400 => x"66c487f5",
  1401 => x"a866c848",
  1402 => x"87cbc004",
  1403 => x"c14866c4",
  1404 => x"58a6c880",
  1405 => x"c887e0c0",
  1406 => x"88c14866",
  1407 => x"c058a6cc",
  1408 => x"c6c187d5",
  1409 => x"c8c005ac",
  1410 => x"4866cc87",
  1411 => x"a6d080c1",
  1412 => x"fcdaff58",
  1413 => x"d04c7087",
  1414 => x"80c14866",
  1415 => x"7458a6d4",
  1416 => x"cbc0029c",
  1417 => x"4866c487",
  1418 => x"a866c8c1",
  1419 => x"87fff204",
  1420 => x"87d4daff",
  1421 => x"c74866c4",
  1422 => x"e5c003a8",
  1423 => x"f4e8c287",
  1424 => x"c478c048",
  1425 => x"91cb4966",
  1426 => x"8166c0c1",
  1427 => x"6a4aa1c4",
  1428 => x"7952c04a",
  1429 => x"c14866c4",
  1430 => x"58a6c880",
  1431 => x"ff04a8c7",
  1432 => x"d0ff87db",
  1433 => x"87fbe08e",
  1434 => x"1e00203a",
  1435 => x"4b711e73",
  1436 => x"87c6029b",
  1437 => x"48f0e8c2",
  1438 => x"1ec778c0",
  1439 => x"bff0e8c2",
  1440 => x"ddc11e49",
  1441 => x"e8c21ed4",
  1442 => x"ee49bfec",
  1443 => x"86cc87f4",
  1444 => x"bfece8c2",
  1445 => x"87f9e949",
  1446 => x"c8029b73",
  1447 => x"d4ddc187",
  1448 => x"e8e5c049",
  1449 => x"fedfff87",
  1450 => x"dac21e87",
  1451 => x"50c048e4",
  1452 => x"bff7dec1",
  1453 => x"c0fbc049",
  1454 => x"2648c087",
  1455 => x"e5c71e4f",
  1456 => x"fe49c187",
  1457 => x"effe87e5",
  1458 => x"987087f1",
  1459 => x"fe87cd02",
  1460 => x"7087eef8",
  1461 => x"87c40298",
  1462 => x"87c24ac1",
  1463 => x"9a724ac0",
  1464 => x"c087ce05",
  1465 => x"cddcc11e",
  1466 => x"eff0c049",
  1467 => x"fe86c487",
  1468 => x"c11ec087",
  1469 => x"c049d8dc",
  1470 => x"c087e1f0",
  1471 => x"87e9fe1e",
  1472 => x"f0c04970",
  1473 => x"dcc387d6",
  1474 => x"268ef887",
  1475 => x"2044534f",
  1476 => x"6c696166",
  1477 => x"002e6465",
  1478 => x"746f6f42",
  1479 => x"2e676e69",
  1480 => x"1e002e2e",
  1481 => x"87c1e8c0",
  1482 => x"87e6f3c0",
  1483 => x"4f2687f6",
  1484 => x"f0e8c21e",
  1485 => x"c278c048",
  1486 => x"c048ece8",
  1487 => x"87fdfd78",
  1488 => x"48c087e1",
  1489 => x"20804f26",
  1490 => x"74697845",
  1491 => x"42208000",
  1492 => x"006b6361",
  1493 => x"000010e9",
  1494 => x"00002a45",
  1495 => x"e9000000",
  1496 => x"63000010",
  1497 => x"0000002a",
  1498 => x"10e90000",
  1499 => x"2a810000",
  1500 => x"00000000",
  1501 => x"0010e900",
  1502 => x"002a9f00",
  1503 => x"00000000",
  1504 => x"000010e9",
  1505 => x"00002abd",
  1506 => x"e9000000",
  1507 => x"db000010",
  1508 => x"0000002a",
  1509 => x"10e90000",
  1510 => x"2af90000",
  1511 => x"00000000",
  1512 => x"0010e900",
  1513 => x"00000000",
  1514 => x"00000000",
  1515 => x"0000117e",
  1516 => x"00000000",
  1517 => x"bb000000",
  1518 => x"42000017",
  1519 => x"20544f4f",
  1520 => x"52202020",
  1521 => x"4c004d4f",
  1522 => x"2064616f",
  1523 => x"1e002e2a",
  1524 => x"c048f0fe",
  1525 => x"7909cd78",
  1526 => x"1e4f2609",
  1527 => x"bff0fe1e",
  1528 => x"2626487e",
  1529 => x"f0fe1e4f",
  1530 => x"2678c148",
  1531 => x"f0fe1e4f",
  1532 => x"2678c048",
  1533 => x"4a711e4f",
  1534 => x"265252c0",
  1535 => x"5b5e0e4f",
  1536 => x"f40e5d5c",
  1537 => x"974d7186",
  1538 => x"a5c17e6d",
  1539 => x"486c974c",
  1540 => x"6e58a6c8",
  1541 => x"a866c448",
  1542 => x"ff87c505",
  1543 => x"87e6c048",
  1544 => x"c287caff",
  1545 => x"6c9749a5",
  1546 => x"4ba3714b",
  1547 => x"974b6b97",
  1548 => x"486e7e6c",
  1549 => x"a6c880c1",
  1550 => x"cc98c758",
  1551 => x"977058a6",
  1552 => x"87e1fe7c",
  1553 => x"8ef44873",
  1554 => x"4c264d26",
  1555 => x"4f264b26",
  1556 => x"5c5b5e0e",
  1557 => x"7186f40e",
  1558 => x"4a66d84c",
  1559 => x"c29affc3",
  1560 => x"6c974ba4",
  1561 => x"49a17349",
  1562 => x"6c975172",
  1563 => x"c1486e7e",
  1564 => x"58a6c880",
  1565 => x"a6cc98c7",
  1566 => x"f4547058",
  1567 => x"87caff8e",
  1568 => x"e8fd1e1e",
  1569 => x"4abfe087",
  1570 => x"c0e0c049",
  1571 => x"87cb0299",
  1572 => x"ecc21e72",
  1573 => x"f7fe49d7",
  1574 => x"fc86c487",
  1575 => x"7e7087fd",
  1576 => x"2687c2fd",
  1577 => x"c21e4f26",
  1578 => x"fd49d7ec",
  1579 => x"e2c187c7",
  1580 => x"dafc49c0",
  1581 => x"87d9c587",
  1582 => x"5e0e4f26",
  1583 => x"0e5d5c5b",
  1584 => x"bff6ecc2",
  1585 => x"cee4c14a",
  1586 => x"724c49bf",
  1587 => x"fc4d71bc",
  1588 => x"4bc087db",
  1589 => x"99d04974",
  1590 => x"7587d502",
  1591 => x"7199d049",
  1592 => x"c11ec01e",
  1593 => x"734ae0ea",
  1594 => x"c0491282",
  1595 => x"86c887e4",
  1596 => x"832d2cc1",
  1597 => x"ff04abc8",
  1598 => x"e8fb87da",
  1599 => x"cee4c187",
  1600 => x"f6ecc248",
  1601 => x"4d2678bf",
  1602 => x"4b264c26",
  1603 => x"00004f26",
  1604 => x"ff1e0000",
  1605 => x"e1c848d0",
  1606 => x"48d4ff78",
  1607 => x"66c478c5",
  1608 => x"c387c302",
  1609 => x"66c878e0",
  1610 => x"ff87c602",
  1611 => x"f0c348d4",
  1612 => x"48d4ff78",
  1613 => x"d0ff7871",
  1614 => x"78e1c848",
  1615 => x"2678e0c0",
  1616 => x"5b5e0e4f",
  1617 => x"4c710e5c",
  1618 => x"49d7ecc2",
  1619 => x"7087eefa",
  1620 => x"aab7c04a",
  1621 => x"87e3c204",
  1622 => x"05aae0c3",
  1623 => x"e8c187c9",
  1624 => x"78c148c4",
  1625 => x"c387d4c2",
  1626 => x"c905aaf0",
  1627 => x"c0e8c187",
  1628 => x"c178c148",
  1629 => x"e8c187f5",
  1630 => x"c702bfc4",
  1631 => x"c24b7287",
  1632 => x"87c2b3c0",
  1633 => x"9c744b72",
  1634 => x"c187d105",
  1635 => x"1ebfc0e8",
  1636 => x"bfc4e8c1",
  1637 => x"fd49721e",
  1638 => x"86c887f8",
  1639 => x"bfc0e8c1",
  1640 => x"87e0c002",
  1641 => x"b7c44973",
  1642 => x"e9c19129",
  1643 => x"4a7381e0",
  1644 => x"92c29acf",
  1645 => x"307248c1",
  1646 => x"baff4a70",
  1647 => x"98694872",
  1648 => x"87db7970",
  1649 => x"b7c44973",
  1650 => x"e9c19129",
  1651 => x"4a7381e0",
  1652 => x"92c29acf",
  1653 => x"307248c3",
  1654 => x"69484a70",
  1655 => x"c17970b0",
  1656 => x"c048c4e8",
  1657 => x"c0e8c178",
  1658 => x"c278c048",
  1659 => x"f849d7ec",
  1660 => x"4a7087cb",
  1661 => x"03aab7c0",
  1662 => x"c087ddfd",
  1663 => x"87c8fc48",
  1664 => x"00000000",
  1665 => x"00000000",
  1666 => x"494a711e",
  1667 => x"2687f2fc",
  1668 => x"4ac01e4f",
  1669 => x"91c44972",
  1670 => x"81e0e9c1",
  1671 => x"82c179c0",
  1672 => x"04aab7d0",
  1673 => x"4f2687ee",
  1674 => x"5c5b5e0e",
  1675 => x"4d710e5d",
  1676 => x"7587faf6",
  1677 => x"2ab7c44a",
  1678 => x"e0e9c192",
  1679 => x"cf4c7582",
  1680 => x"6a94c29c",
  1681 => x"2b744b49",
  1682 => x"48c29bc3",
  1683 => x"4c703074",
  1684 => x"4874bcff",
  1685 => x"7a709871",
  1686 => x"7387caf6",
  1687 => x"87e6fa48",
  1688 => x"00000000",
  1689 => x"00000000",
  1690 => x"00000000",
  1691 => x"00000000",
  1692 => x"00000000",
  1693 => x"00000000",
  1694 => x"00000000",
  1695 => x"00000000",
  1696 => x"00000000",
  1697 => x"00000000",
  1698 => x"00000000",
  1699 => x"00000000",
  1700 => x"00000000",
  1701 => x"00000000",
  1702 => x"00000000",
  1703 => x"00000000",
  1704 => x"25261e16",
  1705 => x"3e3d362e",
  1706 => x"48d0ff1e",
  1707 => x"7178e1c8",
  1708 => x"08d4ff48",
  1709 => x"1e4f2678",
  1710 => x"c848d0ff",
  1711 => x"487178e1",
  1712 => x"7808d4ff",
  1713 => x"ff4866c4",
  1714 => x"267808d4",
  1715 => x"4a711e4f",
  1716 => x"1e4966c4",
  1717 => x"deff4972",
  1718 => x"48d0ff87",
  1719 => x"2678e0c0",
  1720 => x"711e4f26",
  1721 => x"aab7c24a",
  1722 => x"8287c303",
  1723 => x"82ce87c2",
  1724 => x"721e66c4",
  1725 => x"87d5ff49",
  1726 => x"1e4f2626",
  1727 => x"c34ad4ff",
  1728 => x"d0ff7aff",
  1729 => x"78e1c848",
  1730 => x"ecc27ade",
  1731 => x"497abfe1",
  1732 => x"7028c848",
  1733 => x"d048717a",
  1734 => x"717a7028",
  1735 => x"7028d848",
  1736 => x"48d0ff7a",
  1737 => x"2678e0c0",
  1738 => x"5b5e0e4f",
  1739 => x"710e5d5c",
  1740 => x"e1ecc24c",
  1741 => x"744b4dbf",
  1742 => x"9b66d02b",
  1743 => x"66d483c1",
  1744 => x"87c204ab",
  1745 => x"4a744bc0",
  1746 => x"724966d0",
  1747 => x"75b9ff31",
  1748 => x"72487399",
  1749 => x"484a7030",
  1750 => x"ecc2b071",
  1751 => x"dafe58e5",
  1752 => x"264d2687",
  1753 => x"264b264c",
  1754 => x"d0ff1e4f",
  1755 => x"78c9c848",
  1756 => x"d4ff4871",
  1757 => x"4f267808",
  1758 => x"494a711e",
  1759 => x"d0ff87eb",
  1760 => x"2678c848",
  1761 => x"1e731e4f",
  1762 => x"ecc24b71",
  1763 => x"c302bff1",
  1764 => x"87ebc287",
  1765 => x"c848d0ff",
  1766 => x"497378c9",
  1767 => x"ffb1e0c0",
  1768 => x"787148d4",
  1769 => x"48e5ecc2",
  1770 => x"66c878c0",
  1771 => x"c387c502",
  1772 => x"87c249ff",
  1773 => x"ecc249c0",
  1774 => x"66cc59ed",
  1775 => x"c587c602",
  1776 => x"c44ad5d5",
  1777 => x"ffffcf87",
  1778 => x"f1ecc24a",
  1779 => x"f1ecc25a",
  1780 => x"c478c148",
  1781 => x"264d2687",
  1782 => x"264b264c",
  1783 => x"5b5e0e4f",
  1784 => x"710e5d5c",
  1785 => x"edecc24a",
  1786 => x"9a724cbf",
  1787 => x"4987cb02",
  1788 => x"edc191c8",
  1789 => x"83714bfb",
  1790 => x"f1c187c4",
  1791 => x"4dc04bfb",
  1792 => x"99744913",
  1793 => x"bfe9ecc2",
  1794 => x"48d4ffb9",
  1795 => x"b7c17871",
  1796 => x"b7c8852c",
  1797 => x"87e804ad",
  1798 => x"bfe5ecc2",
  1799 => x"c280c848",
  1800 => x"fe58e9ec",
  1801 => x"731e87ef",
  1802 => x"134b711e",
  1803 => x"cb029a4a",
  1804 => x"fe497287",
  1805 => x"4a1387e7",
  1806 => x"87f5059a",
  1807 => x"1e87dafe",
  1808 => x"bfe5ecc2",
  1809 => x"e5ecc249",
  1810 => x"78a1c148",
  1811 => x"a9b7c0c4",
  1812 => x"ff87db03",
  1813 => x"ecc248d4",
  1814 => x"c278bfe9",
  1815 => x"49bfe5ec",
  1816 => x"48e5ecc2",
  1817 => x"c478a1c1",
  1818 => x"04a9b7c0",
  1819 => x"d0ff87e5",
  1820 => x"c278c848",
  1821 => x"c048f1ec",
  1822 => x"004f2678",
  1823 => x"00000000",
  1824 => x"00000000",
  1825 => x"5f5f0000",
  1826 => x"00000000",
  1827 => x"03000303",
  1828 => x"14000003",
  1829 => x"7f147f7f",
  1830 => x"0000147f",
  1831 => x"6b6b2e24",
  1832 => x"4c00123a",
  1833 => x"6c18366a",
  1834 => x"30003256",
  1835 => x"77594f7e",
  1836 => x"0040683a",
  1837 => x"03070400",
  1838 => x"00000000",
  1839 => x"633e1c00",
  1840 => x"00000041",
  1841 => x"3e634100",
  1842 => x"0800001c",
  1843 => x"1c1c3e2a",
  1844 => x"00082a3e",
  1845 => x"3e3e0808",
  1846 => x"00000808",
  1847 => x"60e08000",
  1848 => x"00000000",
  1849 => x"08080808",
  1850 => x"00000808",
  1851 => x"60600000",
  1852 => x"40000000",
  1853 => x"0c183060",
  1854 => x"00010306",
  1855 => x"4d597f3e",
  1856 => x"00003e7f",
  1857 => x"7f7f0604",
  1858 => x"00000000",
  1859 => x"59716342",
  1860 => x"0000464f",
  1861 => x"49496322",
  1862 => x"1800367f",
  1863 => x"7f13161c",
  1864 => x"0000107f",
  1865 => x"45456727",
  1866 => x"0000397d",
  1867 => x"494b7e3c",
  1868 => x"00003079",
  1869 => x"79710101",
  1870 => x"0000070f",
  1871 => x"49497f36",
  1872 => x"0000367f",
  1873 => x"69494f06",
  1874 => x"00001e3f",
  1875 => x"66660000",
  1876 => x"00000000",
  1877 => x"66e68000",
  1878 => x"00000000",
  1879 => x"14140808",
  1880 => x"00002222",
  1881 => x"14141414",
  1882 => x"00001414",
  1883 => x"14142222",
  1884 => x"00000808",
  1885 => x"59510302",
  1886 => x"3e00060f",
  1887 => x"555d417f",
  1888 => x"00001e1f",
  1889 => x"09097f7e",
  1890 => x"00007e7f",
  1891 => x"49497f7f",
  1892 => x"0000367f",
  1893 => x"41633e1c",
  1894 => x"00004141",
  1895 => x"63417f7f",
  1896 => x"00001c3e",
  1897 => x"49497f7f",
  1898 => x"00004141",
  1899 => x"09097f7f",
  1900 => x"00000101",
  1901 => x"49417f3e",
  1902 => x"00007a7b",
  1903 => x"08087f7f",
  1904 => x"00007f7f",
  1905 => x"7f7f4100",
  1906 => x"00000041",
  1907 => x"40406020",
  1908 => x"7f003f7f",
  1909 => x"361c087f",
  1910 => x"00004163",
  1911 => x"40407f7f",
  1912 => x"7f004040",
  1913 => x"060c067f",
  1914 => x"7f007f7f",
  1915 => x"180c067f",
  1916 => x"00007f7f",
  1917 => x"41417f3e",
  1918 => x"00003e7f",
  1919 => x"09097f7f",
  1920 => x"3e00060f",
  1921 => x"7f61417f",
  1922 => x"0000407e",
  1923 => x"19097f7f",
  1924 => x"0000667f",
  1925 => x"594d6f26",
  1926 => x"0000327b",
  1927 => x"7f7f0101",
  1928 => x"00000101",
  1929 => x"40407f3f",
  1930 => x"00003f7f",
  1931 => x"70703f0f",
  1932 => x"7f000f3f",
  1933 => x"3018307f",
  1934 => x"41007f7f",
  1935 => x"1c1c3663",
  1936 => x"01416336",
  1937 => x"7c7c0603",
  1938 => x"61010306",
  1939 => x"474d5971",
  1940 => x"00004143",
  1941 => x"417f7f00",
  1942 => x"01000041",
  1943 => x"180c0603",
  1944 => x"00406030",
  1945 => x"7f414100",
  1946 => x"0800007f",
  1947 => x"0603060c",
  1948 => x"8000080c",
  1949 => x"80808080",
  1950 => x"00008080",
  1951 => x"07030000",
  1952 => x"00000004",
  1953 => x"54547420",
  1954 => x"0000787c",
  1955 => x"44447f7f",
  1956 => x"0000387c",
  1957 => x"44447c38",
  1958 => x"00000044",
  1959 => x"44447c38",
  1960 => x"00007f7f",
  1961 => x"54547c38",
  1962 => x"0000185c",
  1963 => x"057f7e04",
  1964 => x"00000005",
  1965 => x"a4a4bc18",
  1966 => x"00007cfc",
  1967 => x"04047f7f",
  1968 => x"0000787c",
  1969 => x"7d3d0000",
  1970 => x"00000040",
  1971 => x"fd808080",
  1972 => x"0000007d",
  1973 => x"38107f7f",
  1974 => x"0000446c",
  1975 => x"7f3f0000",
  1976 => x"7c000040",
  1977 => x"0c180c7c",
  1978 => x"0000787c",
  1979 => x"04047c7c",
  1980 => x"0000787c",
  1981 => x"44447c38",
  1982 => x"0000387c",
  1983 => x"2424fcfc",
  1984 => x"0000183c",
  1985 => x"24243c18",
  1986 => x"0000fcfc",
  1987 => x"04047c7c",
  1988 => x"0000080c",
  1989 => x"54545c48",
  1990 => x"00002074",
  1991 => x"447f3f04",
  1992 => x"00000044",
  1993 => x"40407c3c",
  1994 => x"00007c7c",
  1995 => x"60603c1c",
  1996 => x"3c001c3c",
  1997 => x"6030607c",
  1998 => x"44003c7c",
  1999 => x"3810386c",
  2000 => x"0000446c",
  2001 => x"60e0bc1c",
  2002 => x"00001c3c",
  2003 => x"5c746444",
  2004 => x"0000444c",
  2005 => x"773e0808",
  2006 => x"00004141",
  2007 => x"7f7f0000",
  2008 => x"00000000",
  2009 => x"3e774141",
  2010 => x"02000808",
  2011 => x"02030101",
  2012 => x"7f000102",
  2013 => x"7f7f7f7f",
  2014 => x"08007f7f",
  2015 => x"3e1c1c08",
  2016 => x"7f7f7f3e",
  2017 => x"1c3e3e7f",
  2018 => x"0008081c",
  2019 => x"7c7c1810",
  2020 => x"00001018",
  2021 => x"7c7c3010",
  2022 => x"10001030",
  2023 => x"78606030",
  2024 => x"4200061e",
  2025 => x"3c183c66",
  2026 => x"78004266",
  2027 => x"c6c26a38",
  2028 => x"6000386c",
  2029 => x"00600000",
  2030 => x"0e006000",
  2031 => x"5d5c5b5e",
  2032 => x"4c711e0e",
  2033 => x"bfc2edc2",
  2034 => x"c04bc04d",
  2035 => x"02ab741e",
  2036 => x"a6c487c7",
  2037 => x"c578c048",
  2038 => x"48a6c487",
  2039 => x"66c478c1",
  2040 => x"ee49731e",
  2041 => x"86c887df",
  2042 => x"ef49e0c0",
  2043 => x"a5c487ef",
  2044 => x"f0496a4a",
  2045 => x"c6f187f0",
  2046 => x"c185cb87",
  2047 => x"abb7c883",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
