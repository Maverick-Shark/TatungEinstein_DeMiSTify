
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"87",x"c7",x"ff",x"04"),
     1 => (x"26",x"4d",x"26",x"26"),
     2 => (x"26",x"4b",x"26",x"4c"),
     3 => (x"4a",x"71",x"1e",x"4f"),
     4 => (x"5a",x"c6",x"ed",x"c2"),
     5 => (x"48",x"c6",x"ed",x"c2"),
     6 => (x"fe",x"49",x"78",x"c7"),
     7 => (x"4f",x"26",x"87",x"dd"),
     8 => (x"71",x"1e",x"73",x"1e"),
     9 => (x"aa",x"b7",x"c0",x"4a"),
    10 => (x"c2",x"87",x"d3",x"03"),
    11 => (x"05",x"bf",x"f1",x"cd"),
    12 => (x"4b",x"c1",x"87",x"c4"),
    13 => (x"4b",x"c0",x"87",x"c2"),
    14 => (x"5b",x"f5",x"cd",x"c2"),
    15 => (x"cd",x"c2",x"87",x"c4"),
    16 => (x"cd",x"c2",x"5a",x"f5"),
    17 => (x"c1",x"4a",x"bf",x"f1"),
    18 => (x"a2",x"c0",x"c1",x"9a"),
    19 => (x"87",x"e8",x"ec",x"49"),
    20 => (x"cd",x"c2",x"48",x"fc"),
    21 => (x"fe",x"78",x"bf",x"f1"),
    22 => (x"71",x"1e",x"87",x"ef"),
    23 => (x"1e",x"66",x"c4",x"4a"),
    24 => (x"fd",x"e9",x"49",x"72"),
    25 => (x"4f",x"26",x"26",x"87"),
    26 => (x"f1",x"cd",x"c2",x"1e"),
    27 => (x"d7",x"e6",x"49",x"bf"),
    28 => (x"fa",x"ec",x"c2",x"87"),
    29 => (x"78",x"bf",x"e8",x"48"),
    30 => (x"48",x"f6",x"ec",x"c2"),
    31 => (x"c2",x"78",x"bf",x"ec"),
    32 => (x"4a",x"bf",x"fa",x"ec"),
    33 => (x"99",x"ff",x"c3",x"49"),
    34 => (x"72",x"2a",x"b7",x"c8"),
    35 => (x"c2",x"b0",x"71",x"48"),
    36 => (x"26",x"58",x"c2",x"ed"),
    37 => (x"5b",x"5e",x"0e",x"4f"),
    38 => (x"71",x"0e",x"5d",x"5c"),
    39 => (x"87",x"c8",x"ff",x"4b"),
    40 => (x"48",x"f5",x"ec",x"c2"),
    41 => (x"49",x"73",x"50",x"c0"),
    42 => (x"70",x"87",x"fd",x"e5"),
    43 => (x"9c",x"c2",x"4c",x"49"),
    44 => (x"cb",x"49",x"ee",x"cb"),
    45 => (x"49",x"70",x"87",x"c3"),
    46 => (x"f5",x"ec",x"c2",x"4d"),
    47 => (x"c1",x"05",x"bf",x"97"),
    48 => (x"66",x"d0",x"87",x"e2"),
    49 => (x"fe",x"ec",x"c2",x"49"),
    50 => (x"d6",x"05",x"99",x"bf"),
    51 => (x"49",x"66",x"d4",x"87"),
    52 => (x"bf",x"f6",x"ec",x"c2"),
    53 => (x"87",x"cb",x"05",x"99"),
    54 => (x"cb",x"e5",x"49",x"73"),
    55 => (x"02",x"98",x"70",x"87"),
    56 => (x"c1",x"87",x"c1",x"c1"),
    57 => (x"87",x"c0",x"fe",x"4c"),
    58 => (x"d8",x"ca",x"49",x"75"),
    59 => (x"02",x"98",x"70",x"87"),
    60 => (x"ec",x"c2",x"87",x"c6"),
    61 => (x"50",x"c1",x"48",x"f5"),
    62 => (x"97",x"f5",x"ec",x"c2"),
    63 => (x"e3",x"c0",x"05",x"bf"),
    64 => (x"fe",x"ec",x"c2",x"87"),
    65 => (x"66",x"d0",x"49",x"bf"),
    66 => (x"d6",x"ff",x"05",x"99"),
    67 => (x"f6",x"ec",x"c2",x"87"),
    68 => (x"66",x"d4",x"49",x"bf"),
    69 => (x"ca",x"ff",x"05",x"99"),
    70 => (x"e4",x"49",x"73",x"87"),
    71 => (x"98",x"70",x"87",x"ca"),
    72 => (x"87",x"ff",x"fe",x"05"),
    73 => (x"dc",x"fb",x"48",x"74"),
    74 => (x"5b",x"5e",x"0e",x"87"),
    75 => (x"f4",x"0e",x"5d",x"5c"),
    76 => (x"4c",x"4d",x"c0",x"86"),
    77 => (x"c4",x"7e",x"bf",x"ec"),
    78 => (x"ed",x"c2",x"48",x"a6"),
    79 => (x"c1",x"78",x"bf",x"c2"),
    80 => (x"c7",x"1e",x"c0",x"1e"),
    81 => (x"87",x"cd",x"fd",x"49"),
    82 => (x"98",x"70",x"86",x"c8"),
    83 => (x"ff",x"87",x"cd",x"02"),
    84 => (x"87",x"cc",x"fb",x"49"),
    85 => (x"e3",x"49",x"da",x"c1"),
    86 => (x"4d",x"c1",x"87",x"ce"),
    87 => (x"97",x"f5",x"ec",x"c2"),
    88 => (x"87",x"c3",x"02",x"bf"),
    89 => (x"c2",x"87",x"fe",x"d4"),
    90 => (x"4b",x"bf",x"fa",x"ec"),
    91 => (x"bf",x"f1",x"cd",x"c2"),
    92 => (x"87",x"e9",x"c0",x"05"),
    93 => (x"e2",x"49",x"fd",x"c3"),
    94 => (x"fa",x"c3",x"87",x"ee"),
    95 => (x"87",x"e8",x"e2",x"49"),
    96 => (x"ff",x"c3",x"49",x"73"),
    97 => (x"c0",x"1e",x"71",x"99"),
    98 => (x"87",x"ce",x"fb",x"49"),
    99 => (x"b7",x"c8",x"49",x"73"),
   100 => (x"c1",x"1e",x"71",x"29"),
   101 => (x"87",x"c2",x"fb",x"49"),
   102 => (x"fa",x"c5",x"86",x"c8"),
   103 => (x"fe",x"ec",x"c2",x"87"),
   104 => (x"02",x"9b",x"4b",x"bf"),
   105 => (x"cd",x"c2",x"87",x"dd"),
   106 => (x"c7",x"49",x"bf",x"ed"),
   107 => (x"98",x"70",x"87",x"d7"),
   108 => (x"c0",x"87",x"c4",x"05"),
   109 => (x"c2",x"87",x"d2",x"4b"),
   110 => (x"fc",x"c6",x"49",x"e0"),
   111 => (x"f1",x"cd",x"c2",x"87"),
   112 => (x"c2",x"87",x"c6",x"58"),
   113 => (x"c0",x"48",x"ed",x"cd"),
   114 => (x"c2",x"49",x"73",x"78"),
   115 => (x"87",x"cd",x"05",x"99"),
   116 => (x"e1",x"49",x"eb",x"c3"),
   117 => (x"49",x"70",x"87",x"d2"),
   118 => (x"c2",x"02",x"99",x"c2"),
   119 => (x"73",x"4c",x"fb",x"87"),
   120 => (x"05",x"99",x"c1",x"49"),
   121 => (x"f4",x"c3",x"87",x"cd"),
   122 => (x"87",x"fc",x"e0",x"49"),
   123 => (x"99",x"c2",x"49",x"70"),
   124 => (x"fa",x"87",x"c2",x"02"),
   125 => (x"c8",x"49",x"73",x"4c"),
   126 => (x"87",x"cd",x"05",x"99"),
   127 => (x"e0",x"49",x"f5",x"c3"),
   128 => (x"49",x"70",x"87",x"e6"),
   129 => (x"d4",x"02",x"99",x"c2"),
   130 => (x"c6",x"ed",x"c2",x"87"),
   131 => (x"87",x"c9",x"02",x"bf"),
   132 => (x"c2",x"88",x"c1",x"48"),
   133 => (x"c2",x"58",x"ca",x"ed"),
   134 => (x"c1",x"4c",x"ff",x"87"),
   135 => (x"c4",x"49",x"73",x"4d"),
   136 => (x"87",x"ce",x"05",x"99"),
   137 => (x"ff",x"49",x"f2",x"c3"),
   138 => (x"70",x"87",x"fd",x"df"),
   139 => (x"02",x"99",x"c2",x"49"),
   140 => (x"ed",x"c2",x"87",x"db"),
   141 => (x"48",x"7e",x"bf",x"c6"),
   142 => (x"03",x"a8",x"b7",x"c7"),
   143 => (x"48",x"6e",x"87",x"cb"),
   144 => (x"ed",x"c2",x"80",x"c1"),
   145 => (x"c2",x"c0",x"58",x"ca"),
   146 => (x"c1",x"4c",x"fe",x"87"),
   147 => (x"49",x"fd",x"c3",x"4d"),
   148 => (x"87",x"d4",x"df",x"ff"),
   149 => (x"99",x"c2",x"49",x"70"),
   150 => (x"c2",x"87",x"d5",x"02"),
   151 => (x"02",x"bf",x"c6",x"ed"),
   152 => (x"c2",x"87",x"c9",x"c0"),
   153 => (x"c0",x"48",x"c6",x"ed"),
   154 => (x"87",x"c2",x"c0",x"78"),
   155 => (x"4d",x"c1",x"4c",x"fd"),
   156 => (x"ff",x"49",x"fa",x"c3"),
   157 => (x"70",x"87",x"f1",x"de"),
   158 => (x"02",x"99",x"c2",x"49"),
   159 => (x"ed",x"c2",x"87",x"d9"),
   160 => (x"c7",x"48",x"bf",x"c6"),
   161 => (x"c0",x"03",x"a8",x"b7"),
   162 => (x"ed",x"c2",x"87",x"c9"),
   163 => (x"78",x"c7",x"48",x"c6"),
   164 => (x"fc",x"87",x"c2",x"c0"),
   165 => (x"c0",x"4d",x"c1",x"4c"),
   166 => (x"c0",x"03",x"ac",x"b7"),
   167 => (x"66",x"c4",x"87",x"d1"),
   168 => (x"82",x"d8",x"c1",x"4a"),
   169 => (x"c6",x"c0",x"02",x"6a"),
   170 => (x"74",x"4b",x"6a",x"87"),
   171 => (x"c0",x"0f",x"73",x"49"),
   172 => (x"1e",x"f0",x"c3",x"1e"),
   173 => (x"f7",x"49",x"da",x"c1"),
   174 => (x"86",x"c8",x"87",x"db"),
   175 => (x"c0",x"02",x"98",x"70"),
   176 => (x"a6",x"c8",x"87",x"e2"),
   177 => (x"c6",x"ed",x"c2",x"48"),
   178 => (x"66",x"c8",x"78",x"bf"),
   179 => (x"c4",x"91",x"cb",x"49"),
   180 => (x"80",x"71",x"48",x"66"),
   181 => (x"bf",x"6e",x"7e",x"70"),
   182 => (x"87",x"c8",x"c0",x"02"),
   183 => (x"c8",x"4b",x"bf",x"6e"),
   184 => (x"0f",x"73",x"49",x"66"),
   185 => (x"c0",x"02",x"9d",x"75"),
   186 => (x"ed",x"c2",x"87",x"c8"),
   187 => (x"f3",x"49",x"bf",x"c6"),
   188 => (x"cd",x"c2",x"87",x"c9"),
   189 => (x"c0",x"02",x"bf",x"f5"),
   190 => (x"c2",x"49",x"87",x"dd"),
   191 => (x"98",x"70",x"87",x"c7"),
   192 => (x"87",x"d3",x"c0",x"02"),
   193 => (x"bf",x"c6",x"ed",x"c2"),
   194 => (x"87",x"ef",x"f2",x"49"),
   195 => (x"cf",x"f4",x"49",x"c0"),
   196 => (x"f5",x"cd",x"c2",x"87"),
   197 => (x"f4",x"78",x"c0",x"48"),
   198 => (x"87",x"e9",x"f3",x"8e"),
   199 => (x"5c",x"5b",x"5e",x"0e"),
   200 => (x"71",x"1e",x"0e",x"5d"),
   201 => (x"c2",x"ed",x"c2",x"4c"),
   202 => (x"cd",x"c1",x"49",x"bf"),
   203 => (x"d1",x"c1",x"4d",x"a1"),
   204 => (x"74",x"7e",x"69",x"81"),
   205 => (x"87",x"cf",x"02",x"9c"),
   206 => (x"74",x"4b",x"a5",x"c4"),
   207 => (x"c2",x"ed",x"c2",x"7b"),
   208 => (x"c8",x"f3",x"49",x"bf"),
   209 => (x"74",x"7b",x"6e",x"87"),
   210 => (x"87",x"c4",x"05",x"9c"),
   211 => (x"87",x"c2",x"4b",x"c0"),
   212 => (x"49",x"73",x"4b",x"c1"),
   213 => (x"d4",x"87",x"c9",x"f3"),
   214 => (x"87",x"c7",x"02",x"66"),
   215 => (x"70",x"87",x"da",x"49"),
   216 => (x"c0",x"87",x"c2",x"4a"),
   217 => (x"f9",x"cd",x"c2",x"4a"),
   218 => (x"d8",x"f2",x"26",x"5a"),
   219 => (x"00",x"00",x"00",x"87"),
   220 => (x"00",x"00",x"00",x"00"),
   221 => (x"00",x"00",x"00",x"00"),
   222 => (x"4a",x"71",x"1e",x"00"),
   223 => (x"49",x"bf",x"c8",x"ff"),
   224 => (x"26",x"48",x"a1",x"72"),
   225 => (x"c8",x"ff",x"1e",x"4f"),
   226 => (x"c0",x"fe",x"89",x"bf"),
   227 => (x"c0",x"c0",x"c0",x"c0"),
   228 => (x"87",x"c4",x"01",x"a9"),
   229 => (x"87",x"c2",x"4a",x"c0"),
   230 => (x"48",x"72",x"4a",x"c1"),
   231 => (x"5e",x"0e",x"4f",x"26"),
   232 => (x"0e",x"5d",x"5c",x"5b"),
   233 => (x"d4",x"ff",x"4b",x"71"),
   234 => (x"48",x"66",x"d0",x"4c"),
   235 => (x"49",x"d6",x"78",x"c0"),
   236 => (x"87",x"f4",x"db",x"ff"),
   237 => (x"6c",x"7c",x"ff",x"c3"),
   238 => (x"99",x"ff",x"c3",x"49"),
   239 => (x"c3",x"49",x"4d",x"71"),
   240 => (x"e0",x"c1",x"99",x"f0"),
   241 => (x"87",x"cb",x"05",x"a9"),
   242 => (x"6c",x"7c",x"ff",x"c3"),
   243 => (x"d0",x"98",x"c3",x"48"),
   244 => (x"c3",x"78",x"08",x"66"),
   245 => (x"4a",x"6c",x"7c",x"ff"),
   246 => (x"c3",x"31",x"c8",x"49"),
   247 => (x"4a",x"6c",x"7c",x"ff"),
   248 => (x"49",x"72",x"b2",x"71"),
   249 => (x"ff",x"c3",x"31",x"c8"),
   250 => (x"71",x"4a",x"6c",x"7c"),
   251 => (x"c8",x"49",x"72",x"b2"),
   252 => (x"7c",x"ff",x"c3",x"31"),
   253 => (x"b2",x"71",x"4a",x"6c"),
   254 => (x"c0",x"48",x"d0",x"ff"),
   255 => (x"9b",x"73",x"78",x"e0"),
   256 => (x"72",x"87",x"c2",x"02"),
   257 => (x"26",x"48",x"75",x"7b"),
   258 => (x"26",x"4c",x"26",x"4d"),
   259 => (x"1e",x"4f",x"26",x"4b"),
   260 => (x"5e",x"0e",x"4f",x"26"),
   261 => (x"f8",x"0e",x"5c",x"5b"),
   262 => (x"c8",x"1e",x"76",x"86"),
   263 => (x"fd",x"fd",x"49",x"a6"),
   264 => (x"70",x"86",x"c4",x"87"),
   265 => (x"c0",x"48",x"6e",x"4b"),
   266 => (x"c6",x"c3",x"01",x"a8"),
   267 => (x"c3",x"4a",x"73",x"87"),
   268 => (x"d0",x"c1",x"9a",x"f0"),
   269 => (x"87",x"c7",x"02",x"aa"),
   270 => (x"05",x"aa",x"e0",x"c1"),
   271 => (x"73",x"87",x"f4",x"c2"),
   272 => (x"02",x"99",x"c8",x"49"),
   273 => (x"c6",x"ff",x"87",x"c3"),
   274 => (x"c3",x"4c",x"73",x"87"),
   275 => (x"05",x"ac",x"c2",x"9c"),
   276 => (x"c4",x"87",x"cd",x"c1"),
   277 => (x"31",x"c9",x"49",x"66"),
   278 => (x"66",x"c4",x"1e",x"71"),
   279 => (x"c2",x"92",x"d4",x"4a"),
   280 => (x"72",x"49",x"ca",x"ed"),
   281 => (x"c6",x"d5",x"fe",x"81"),
   282 => (x"49",x"66",x"c4",x"87"),
   283 => (x"49",x"e3",x"c0",x"1e"),
   284 => (x"87",x"d9",x"d9",x"ff"),
   285 => (x"d8",x"ff",x"49",x"d8"),
   286 => (x"c0",x"c8",x"87",x"ee"),
   287 => (x"fa",x"db",x"c2",x"1e"),
   288 => (x"d6",x"f1",x"fd",x"49"),
   289 => (x"48",x"d0",x"ff",x"87"),
   290 => (x"c2",x"78",x"e0",x"c0"),
   291 => (x"d0",x"1e",x"fa",x"db"),
   292 => (x"92",x"d4",x"4a",x"66"),
   293 => (x"49",x"ca",x"ed",x"c2"),
   294 => (x"d3",x"fe",x"81",x"72"),
   295 => (x"86",x"d0",x"87",x"ce"),
   296 => (x"c1",x"05",x"ac",x"c1"),
   297 => (x"66",x"c4",x"87",x"cd"),
   298 => (x"71",x"31",x"c9",x"49"),
   299 => (x"4a",x"66",x"c4",x"1e"),
   300 => (x"ed",x"c2",x"92",x"d4"),
   301 => (x"81",x"72",x"49",x"ca"),
   302 => (x"87",x"f3",x"d3",x"fe"),
   303 => (x"1e",x"fa",x"db",x"c2"),
   304 => (x"d4",x"4a",x"66",x"c8"),
   305 => (x"ca",x"ed",x"c2",x"92"),
   306 => (x"fe",x"81",x"72",x"49"),
   307 => (x"c8",x"87",x"da",x"d1"),
   308 => (x"c0",x"1e",x"49",x"66"),
   309 => (x"d7",x"ff",x"49",x"e3"),
   310 => (x"49",x"d7",x"87",x"f3"),
   311 => (x"87",x"c8",x"d7",x"ff"),
   312 => (x"c2",x"1e",x"c0",x"c8"),
   313 => (x"fd",x"49",x"fa",x"db"),
   314 => (x"d0",x"87",x"da",x"ef"),
   315 => (x"48",x"d0",x"ff",x"86"),
   316 => (x"f8",x"78",x"e0",x"c0"),
   317 => (x"87",x"d1",x"fc",x"8e"),
   318 => (x"5c",x"5b",x"5e",x"0e"),
   319 => (x"71",x"1e",x"0e",x"5d"),
   320 => (x"4c",x"d4",x"ff",x"4d"),
   321 => (x"48",x"7e",x"66",x"d4"),
   322 => (x"06",x"a8",x"b7",x"c3"),
   323 => (x"48",x"c0",x"87",x"c5"),
   324 => (x"75",x"87",x"e2",x"c1"),
   325 => (x"e7",x"e1",x"fe",x"49"),
   326 => (x"c4",x"1e",x"75",x"87"),
   327 => (x"93",x"d4",x"4b",x"66"),
   328 => (x"83",x"ca",x"ed",x"c2"),
   329 => (x"cc",x"fe",x"49",x"73"),
   330 => (x"83",x"c8",x"87",x"e3"),
   331 => (x"d0",x"ff",x"4b",x"6b"),
   332 => (x"78",x"e1",x"c8",x"48"),
   333 => (x"49",x"73",x"7c",x"dd"),
   334 => (x"71",x"99",x"ff",x"c3"),
   335 => (x"c8",x"49",x"73",x"7c"),
   336 => (x"ff",x"c3",x"29",x"b7"),
   337 => (x"73",x"7c",x"71",x"99"),
   338 => (x"29",x"b7",x"d0",x"49"),
   339 => (x"71",x"99",x"ff",x"c3"),
   340 => (x"d8",x"49",x"73",x"7c"),
   341 => (x"7c",x"71",x"29",x"b7"),
   342 => (x"7c",x"7c",x"7c",x"c0"),
   343 => (x"7c",x"7c",x"7c",x"7c"),
   344 => (x"7c",x"7c",x"7c",x"7c"),
   345 => (x"78",x"e0",x"c0",x"7c"),
   346 => (x"dc",x"1e",x"66",x"c4"),
   347 => (x"dc",x"d5",x"ff",x"49"),
   348 => (x"73",x"86",x"c8",x"87"),
   349 => (x"ce",x"fa",x"26",x"48"),
   350 => (x"5b",x"5e",x"0e",x"87"),
   351 => (x"1e",x"0e",x"5d",x"5c"),
   352 => (x"d4",x"ff",x"7e",x"71"),
   353 => (x"c2",x"1e",x"6e",x"4b"),
   354 => (x"fe",x"49",x"de",x"ed"),
   355 => (x"c4",x"87",x"fe",x"ca"),
   356 => (x"9d",x"4d",x"70",x"86"),
   357 => (x"87",x"c3",x"c3",x"02"),
   358 => (x"bf",x"e6",x"ed",x"c2"),
   359 => (x"fe",x"49",x"6e",x"4c"),
   360 => (x"ff",x"87",x"dd",x"df"),
   361 => (x"c5",x"c8",x"48",x"d0"),
   362 => (x"7b",x"d6",x"c1",x"78"),
   363 => (x"7b",x"15",x"4a",x"c0"),
   364 => (x"e0",x"c0",x"82",x"c1"),
   365 => (x"f5",x"04",x"aa",x"b7"),
   366 => (x"48",x"d0",x"ff",x"87"),
   367 => (x"c5",x"c8",x"78",x"c4"),
   368 => (x"7b",x"d3",x"c1",x"78"),
   369 => (x"78",x"c4",x"7b",x"c1"),
   370 => (x"c1",x"02",x"9c",x"74"),
   371 => (x"db",x"c2",x"87",x"fc"),
   372 => (x"c0",x"c8",x"7e",x"fa"),
   373 => (x"b7",x"c0",x"8c",x"4d"),
   374 => (x"87",x"c6",x"03",x"ac"),
   375 => (x"4d",x"a4",x"c0",x"c8"),
   376 => (x"e8",x"c2",x"4c",x"c0"),
   377 => (x"49",x"bf",x"97",x"eb"),
   378 => (x"d2",x"02",x"99",x"d0"),
   379 => (x"c2",x"1e",x"c0",x"87"),
   380 => (x"fe",x"49",x"de",x"ed"),
   381 => (x"c4",x"87",x"f2",x"cc"),
   382 => (x"4a",x"49",x"70",x"86"),
   383 => (x"c2",x"87",x"ef",x"c0"),
   384 => (x"c2",x"1e",x"fa",x"db"),
   385 => (x"fe",x"49",x"de",x"ed"),
   386 => (x"c4",x"87",x"de",x"cc"),
   387 => (x"4a",x"49",x"70",x"86"),
   388 => (x"c8",x"48",x"d0",x"ff"),
   389 => (x"d4",x"c1",x"78",x"c5"),
   390 => (x"bf",x"97",x"6e",x"7b"),
   391 => (x"c1",x"48",x"6e",x"7b"),
   392 => (x"c1",x"7e",x"70",x"80"),
   393 => (x"f0",x"ff",x"05",x"8d"),
   394 => (x"48",x"d0",x"ff",x"87"),
   395 => (x"9a",x"72",x"78",x"c4"),
   396 => (x"c0",x"87",x"c5",x"05"),
   397 => (x"87",x"e5",x"c0",x"48"),
   398 => (x"ed",x"c2",x"1e",x"c1"),
   399 => (x"ca",x"fe",x"49",x"de"),
   400 => (x"86",x"c4",x"87",x"c6"),
   401 => (x"fe",x"05",x"9c",x"74"),
   402 => (x"d0",x"ff",x"87",x"c4"),
   403 => (x"78",x"c5",x"c8",x"48"),
   404 => (x"c0",x"7b",x"d3",x"c1"),
   405 => (x"c1",x"78",x"c4",x"7b"),
   406 => (x"c0",x"87",x"c2",x"48"),
   407 => (x"4d",x"26",x"26",x"48"),
   408 => (x"4b",x"26",x"4c",x"26"),
   409 => (x"5e",x"0e",x"4f",x"26"),
   410 => (x"71",x"0e",x"5c",x"5b"),
   411 => (x"02",x"66",x"cc",x"4b"),
   412 => (x"c0",x"4c",x"87",x"d8"),
   413 => (x"d8",x"02",x"8c",x"f0"),
   414 => (x"c1",x"4a",x"74",x"87"),
   415 => (x"87",x"d1",x"02",x"8a"),
   416 => (x"87",x"cd",x"02",x"8a"),
   417 => (x"87",x"c9",x"02",x"8a"),
   418 => (x"49",x"73",x"87",x"d7"),
   419 => (x"d0",x"87",x"ea",x"fb"),
   420 => (x"c0",x"1e",x"74",x"87"),
   421 => (x"87",x"e0",x"f9",x"49"),
   422 => (x"49",x"73",x"1e",x"74"),
   423 => (x"c8",x"87",x"d9",x"f9"),
   424 => (x"87",x"fc",x"fe",x"86"),
   425 => (x"db",x"c2",x"1e",x"00"),
   426 => (x"c1",x"49",x"bf",x"ce"),
   427 => (x"d2",x"db",x"c2",x"b9"),
   428 => (x"48",x"d4",x"ff",x"59"),
   429 => (x"ff",x"78",x"ff",x"c3"),
   430 => (x"e1",x"c8",x"48",x"d0"),
   431 => (x"48",x"d4",x"ff",x"78"),
   432 => (x"31",x"c4",x"78",x"c1"),
   433 => (x"d0",x"ff",x"78",x"71"),
   434 => (x"78",x"e0",x"c0",x"48"),
   435 => (x"00",x"00",x"4f",x"26"),
   436 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

