library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"87c7ff04",
     1 => x"264d2626",
     2 => x"264b264c",
     3 => x"4a711e4f",
     4 => x"5ac6edc2",
     5 => x"48c6edc2",
     6 => x"fe4978c7",
     7 => x"4f2687dd",
     8 => x"711e731e",
     9 => x"aab7c04a",
    10 => x"c287d303",
    11 => x"05bff1cd",
    12 => x"4bc187c4",
    13 => x"4bc087c2",
    14 => x"5bf5cdc2",
    15 => x"cdc287c4",
    16 => x"cdc25af5",
    17 => x"c14abff1",
    18 => x"a2c0c19a",
    19 => x"87e8ec49",
    20 => x"cdc248fc",
    21 => x"fe78bff1",
    22 => x"711e87ef",
    23 => x"1e66c44a",
    24 => x"fde94972",
    25 => x"4f262687",
    26 => x"f1cdc21e",
    27 => x"d7e649bf",
    28 => x"faecc287",
    29 => x"78bfe848",
    30 => x"48f6ecc2",
    31 => x"c278bfec",
    32 => x"4abffaec",
    33 => x"99ffc349",
    34 => x"722ab7c8",
    35 => x"c2b07148",
    36 => x"2658c2ed",
    37 => x"5b5e0e4f",
    38 => x"710e5d5c",
    39 => x"87c8ff4b",
    40 => x"48f5ecc2",
    41 => x"497350c0",
    42 => x"7087fde5",
    43 => x"9cc24c49",
    44 => x"cb49eecb",
    45 => x"497087c3",
    46 => x"f5ecc24d",
    47 => x"c105bf97",
    48 => x"66d087e2",
    49 => x"feecc249",
    50 => x"d60599bf",
    51 => x"4966d487",
    52 => x"bff6ecc2",
    53 => x"87cb0599",
    54 => x"cbe54973",
    55 => x"02987087",
    56 => x"c187c1c1",
    57 => x"87c0fe4c",
    58 => x"d8ca4975",
    59 => x"02987087",
    60 => x"ecc287c6",
    61 => x"50c148f5",
    62 => x"97f5ecc2",
    63 => x"e3c005bf",
    64 => x"feecc287",
    65 => x"66d049bf",
    66 => x"d6ff0599",
    67 => x"f6ecc287",
    68 => x"66d449bf",
    69 => x"caff0599",
    70 => x"e4497387",
    71 => x"987087ca",
    72 => x"87fffe05",
    73 => x"dcfb4874",
    74 => x"5b5e0e87",
    75 => x"f40e5d5c",
    76 => x"4c4dc086",
    77 => x"c47ebfec",
    78 => x"edc248a6",
    79 => x"c178bfc2",
    80 => x"c71ec01e",
    81 => x"87cdfd49",
    82 => x"987086c8",
    83 => x"ff87cd02",
    84 => x"87ccfb49",
    85 => x"e349dac1",
    86 => x"4dc187ce",
    87 => x"97f5ecc2",
    88 => x"87c302bf",
    89 => x"c287fed4",
    90 => x"4bbffaec",
    91 => x"bff1cdc2",
    92 => x"87e9c005",
    93 => x"e249fdc3",
    94 => x"fac387ee",
    95 => x"87e8e249",
    96 => x"ffc34973",
    97 => x"c01e7199",
    98 => x"87cefb49",
    99 => x"b7c84973",
   100 => x"c11e7129",
   101 => x"87c2fb49",
   102 => x"fac586c8",
   103 => x"feecc287",
   104 => x"029b4bbf",
   105 => x"cdc287dd",
   106 => x"c749bfed",
   107 => x"987087d7",
   108 => x"c087c405",
   109 => x"c287d24b",
   110 => x"fcc649e0",
   111 => x"f1cdc287",
   112 => x"c287c658",
   113 => x"c048edcd",
   114 => x"c2497378",
   115 => x"87cd0599",
   116 => x"e149ebc3",
   117 => x"497087d2",
   118 => x"c20299c2",
   119 => x"734cfb87",
   120 => x"0599c149",
   121 => x"f4c387cd",
   122 => x"87fce049",
   123 => x"99c24970",
   124 => x"fa87c202",
   125 => x"c849734c",
   126 => x"87cd0599",
   127 => x"e049f5c3",
   128 => x"497087e6",
   129 => x"d40299c2",
   130 => x"c6edc287",
   131 => x"87c902bf",
   132 => x"c288c148",
   133 => x"c258caed",
   134 => x"c14cff87",
   135 => x"c449734d",
   136 => x"87ce0599",
   137 => x"ff49f2c3",
   138 => x"7087fddf",
   139 => x"0299c249",
   140 => x"edc287db",
   141 => x"487ebfc6",
   142 => x"03a8b7c7",
   143 => x"486e87cb",
   144 => x"edc280c1",
   145 => x"c2c058ca",
   146 => x"c14cfe87",
   147 => x"49fdc34d",
   148 => x"87d4dfff",
   149 => x"99c24970",
   150 => x"c287d502",
   151 => x"02bfc6ed",
   152 => x"c287c9c0",
   153 => x"c048c6ed",
   154 => x"87c2c078",
   155 => x"4dc14cfd",
   156 => x"ff49fac3",
   157 => x"7087f1de",
   158 => x"0299c249",
   159 => x"edc287d9",
   160 => x"c748bfc6",
   161 => x"c003a8b7",
   162 => x"edc287c9",
   163 => x"78c748c6",
   164 => x"fc87c2c0",
   165 => x"c04dc14c",
   166 => x"c003acb7",
   167 => x"66c487d1",
   168 => x"82d8c14a",
   169 => x"c6c0026a",
   170 => x"744b6a87",
   171 => x"c00f7349",
   172 => x"1ef0c31e",
   173 => x"f749dac1",
   174 => x"86c887db",
   175 => x"c0029870",
   176 => x"a6c887e2",
   177 => x"c6edc248",
   178 => x"66c878bf",
   179 => x"c491cb49",
   180 => x"80714866",
   181 => x"bf6e7e70",
   182 => x"87c8c002",
   183 => x"c84bbf6e",
   184 => x"0f734966",
   185 => x"c0029d75",
   186 => x"edc287c8",
   187 => x"f349bfc6",
   188 => x"cdc287c9",
   189 => x"c002bff5",
   190 => x"c24987dd",
   191 => x"987087c7",
   192 => x"87d3c002",
   193 => x"bfc6edc2",
   194 => x"87eff249",
   195 => x"cff449c0",
   196 => x"f5cdc287",
   197 => x"f478c048",
   198 => x"87e9f38e",
   199 => x"5c5b5e0e",
   200 => x"711e0e5d",
   201 => x"c2edc24c",
   202 => x"cdc149bf",
   203 => x"d1c14da1",
   204 => x"747e6981",
   205 => x"87cf029c",
   206 => x"744ba5c4",
   207 => x"c2edc27b",
   208 => x"c8f349bf",
   209 => x"747b6e87",
   210 => x"87c4059c",
   211 => x"87c24bc0",
   212 => x"49734bc1",
   213 => x"d487c9f3",
   214 => x"87c70266",
   215 => x"7087da49",
   216 => x"c087c24a",
   217 => x"f9cdc24a",
   218 => x"d8f2265a",
   219 => x"00000087",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"4a711e00",
   223 => x"49bfc8ff",
   224 => x"2648a172",
   225 => x"c8ff1e4f",
   226 => x"c0fe89bf",
   227 => x"c0c0c0c0",
   228 => x"87c401a9",
   229 => x"87c24ac0",
   230 => x"48724ac1",
   231 => x"5e0e4f26",
   232 => x"0e5d5c5b",
   233 => x"d4ff4b71",
   234 => x"4866d04c",
   235 => x"49d678c0",
   236 => x"87f4dbff",
   237 => x"6c7cffc3",
   238 => x"99ffc349",
   239 => x"c3494d71",
   240 => x"e0c199f0",
   241 => x"87cb05a9",
   242 => x"6c7cffc3",
   243 => x"d098c348",
   244 => x"c3780866",
   245 => x"4a6c7cff",
   246 => x"c331c849",
   247 => x"4a6c7cff",
   248 => x"4972b271",
   249 => x"ffc331c8",
   250 => x"714a6c7c",
   251 => x"c84972b2",
   252 => x"7cffc331",
   253 => x"b2714a6c",
   254 => x"c048d0ff",
   255 => x"9b7378e0",
   256 => x"7287c202",
   257 => x"2648757b",
   258 => x"264c264d",
   259 => x"1e4f264b",
   260 => x"5e0e4f26",
   261 => x"f80e5c5b",
   262 => x"c81e7686",
   263 => x"fdfd49a6",
   264 => x"7086c487",
   265 => x"c0486e4b",
   266 => x"c6c301a8",
   267 => x"c34a7387",
   268 => x"d0c19af0",
   269 => x"87c702aa",
   270 => x"05aae0c1",
   271 => x"7387f4c2",
   272 => x"0299c849",
   273 => x"c6ff87c3",
   274 => x"c34c7387",
   275 => x"05acc29c",
   276 => x"c487cdc1",
   277 => x"31c94966",
   278 => x"66c41e71",
   279 => x"c292d44a",
   280 => x"7249caed",
   281 => x"c6d5fe81",
   282 => x"4966c487",
   283 => x"49e3c01e",
   284 => x"87d9d9ff",
   285 => x"d8ff49d8",
   286 => x"c0c887ee",
   287 => x"fadbc21e",
   288 => x"d6f1fd49",
   289 => x"48d0ff87",
   290 => x"c278e0c0",
   291 => x"d01efadb",
   292 => x"92d44a66",
   293 => x"49caedc2",
   294 => x"d3fe8172",
   295 => x"86d087ce",
   296 => x"c105acc1",
   297 => x"66c487cd",
   298 => x"7131c949",
   299 => x"4a66c41e",
   300 => x"edc292d4",
   301 => x"817249ca",
   302 => x"87f3d3fe",
   303 => x"1efadbc2",
   304 => x"d44a66c8",
   305 => x"caedc292",
   306 => x"fe817249",
   307 => x"c887dad1",
   308 => x"c01e4966",
   309 => x"d7ff49e3",
   310 => x"49d787f3",
   311 => x"87c8d7ff",
   312 => x"c21ec0c8",
   313 => x"fd49fadb",
   314 => x"d087daef",
   315 => x"48d0ff86",
   316 => x"f878e0c0",
   317 => x"87d1fc8e",
   318 => x"5c5b5e0e",
   319 => x"711e0e5d",
   320 => x"4cd4ff4d",
   321 => x"487e66d4",
   322 => x"06a8b7c3",
   323 => x"48c087c5",
   324 => x"7587e2c1",
   325 => x"e7e1fe49",
   326 => x"c41e7587",
   327 => x"93d44b66",
   328 => x"83caedc2",
   329 => x"ccfe4973",
   330 => x"83c887e3",
   331 => x"d0ff4b6b",
   332 => x"78e1c848",
   333 => x"49737cdd",
   334 => x"7199ffc3",
   335 => x"c849737c",
   336 => x"ffc329b7",
   337 => x"737c7199",
   338 => x"29b7d049",
   339 => x"7199ffc3",
   340 => x"d849737c",
   341 => x"7c7129b7",
   342 => x"7c7c7cc0",
   343 => x"7c7c7c7c",
   344 => x"7c7c7c7c",
   345 => x"78e0c07c",
   346 => x"dc1e66c4",
   347 => x"dcd5ff49",
   348 => x"7386c887",
   349 => x"cefa2648",
   350 => x"5b5e0e87",
   351 => x"1e0e5d5c",
   352 => x"d4ff7e71",
   353 => x"c21e6e4b",
   354 => x"fe49deed",
   355 => x"c487feca",
   356 => x"9d4d7086",
   357 => x"87c3c302",
   358 => x"bfe6edc2",
   359 => x"fe496e4c",
   360 => x"ff87dddf",
   361 => x"c5c848d0",
   362 => x"7bd6c178",
   363 => x"7b154ac0",
   364 => x"e0c082c1",
   365 => x"f504aab7",
   366 => x"48d0ff87",
   367 => x"c5c878c4",
   368 => x"7bd3c178",
   369 => x"78c47bc1",
   370 => x"c1029c74",
   371 => x"dbc287fc",
   372 => x"c0c87efa",
   373 => x"b7c08c4d",
   374 => x"87c603ac",
   375 => x"4da4c0c8",
   376 => x"e8c24cc0",
   377 => x"49bf97eb",
   378 => x"d20299d0",
   379 => x"c21ec087",
   380 => x"fe49deed",
   381 => x"c487f2cc",
   382 => x"4a497086",
   383 => x"c287efc0",
   384 => x"c21efadb",
   385 => x"fe49deed",
   386 => x"c487decc",
   387 => x"4a497086",
   388 => x"c848d0ff",
   389 => x"d4c178c5",
   390 => x"bf976e7b",
   391 => x"c1486e7b",
   392 => x"c17e7080",
   393 => x"f0ff058d",
   394 => x"48d0ff87",
   395 => x"9a7278c4",
   396 => x"c087c505",
   397 => x"87e5c048",
   398 => x"edc21ec1",
   399 => x"cafe49de",
   400 => x"86c487c6",
   401 => x"fe059c74",
   402 => x"d0ff87c4",
   403 => x"78c5c848",
   404 => x"c07bd3c1",
   405 => x"c178c47b",
   406 => x"c087c248",
   407 => x"4d262648",
   408 => x"4b264c26",
   409 => x"5e0e4f26",
   410 => x"710e5c5b",
   411 => x"0266cc4b",
   412 => x"c04c87d8",
   413 => x"d8028cf0",
   414 => x"c14a7487",
   415 => x"87d1028a",
   416 => x"87cd028a",
   417 => x"87c9028a",
   418 => x"497387d7",
   419 => x"d087eafb",
   420 => x"c01e7487",
   421 => x"87e0f949",
   422 => x"49731e74",
   423 => x"c887d9f9",
   424 => x"87fcfe86",
   425 => x"dbc21e00",
   426 => x"c149bfce",
   427 => x"d2dbc2b9",
   428 => x"48d4ff59",
   429 => x"ff78ffc3",
   430 => x"e1c848d0",
   431 => x"48d4ff78",
   432 => x"31c478c1",
   433 => x"d0ff7871",
   434 => x"78e0c048",
   435 => x"00004f26",
   436 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
